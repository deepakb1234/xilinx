always@(reset)
begin
reg_space[1024] = 8'h00;
reg_space[1025] = 8'h00;
reg_space[1026] = 8'h00;
reg_space[1027] = 8'h00;
reg_space[1028] = 8'h00;
reg_space[1029] = 8'h00;
reg_space[1030] = 8'h00;
reg_space[1031] = 8'h00;
reg_space[1032] = 8'h00;
reg_space[1033] = 8'h00;
reg_space[1034] = 8'h00;
reg_space[1035] = 8'h00;
reg_space[1036] = 8'h00;
reg_space[1037] = 8'h00;
reg_space[1038] = 8'h00;
reg_space[1039] = 8'h00;
reg_space[1040] = 8'h00;
reg_space[1041] = 8'h00;
reg_space[1042] = 8'h00;
reg_space[1043] = 8'h00;
reg_space[1044] = 8'h00;
reg_space[1045] = 8'h00;
reg_space[1046] = 8'h00;
reg_space[1047] = 8'h00;
reg_space[1048] = 8'h00;
reg_space[1049] = 8'h00;
reg_space[1050] = 8'h00;
reg_space[1051] = 8'h00;
reg_space[1052] = 8'h00;
reg_space[1053] = 8'h00;
reg_space[1054] = 8'h00;
reg_space[1055] = 8'h00;
reg_space[1056] = 8'h00;
reg_space[1057] = 8'h00;
reg_space[1058] = 8'h00;
reg_space[1059] = 8'h00;
reg_space[1060] = 8'h00;
reg_space[1061] = 8'h00;
reg_space[1062] = 8'h00;
reg_space[1063] = 8'h00;
reg_space[1064] = 8'h00;
reg_space[1065] = 8'h00;
reg_space[1066] = 8'h00;
reg_space[1067] = 8'h00;
reg_space[1068] = 8'h00;
reg_space[1069] = 8'h00;
reg_space[1070] = 8'h00;
reg_space[1071] = 8'h00;
reg_space[1072] = 8'h00;
reg_space[1073] = 8'h00;
reg_space[1074] = 8'h00;
reg_space[1075] = 8'h00;
reg_space[1076] = 8'h00;
reg_space[1077] = 8'h00;
reg_space[1078] = 8'h00;
reg_space[1079] = 8'h00;
reg_space[1080] = 8'h00;
reg_space[1081] = 8'h00;
reg_space[1082] = 8'h00;
reg_space[1083] = 8'h00;
reg_space[1084] = 8'h00;
reg_space[1085] = 8'h00;
reg_space[1086] = 8'h00;
reg_space[1087] = 8'h00;
reg_space[1088] = 8'h00;
reg_space[1089] = 8'h00;
reg_space[1090] = 8'h00;
reg_space[1091] = 8'h00;
reg_space[1092] = 8'h00;
reg_space[1093] = 8'h00;
reg_space[1094] = 8'h00;
reg_space[1095] = 8'h00;
reg_space[1096] = 8'h00;
reg_space[1097] = 8'h00;
reg_space[1098] = 8'h00;
reg_space[1099] = 8'h00;
reg_space[1100] = 8'h00;
reg_space[1101] = 8'h00;
reg_space[1102] = 8'h00;
reg_space[1103] = 8'h00;
reg_space[1104] = 8'h00;
reg_space[1105] = 8'h00;
reg_space[1106] = 8'h00;
reg_space[1107] = 8'h00;
reg_space[1108] = 8'h00;
reg_space[1109] = 8'h00;
reg_space[1110] = 8'h00;
reg_space[1111] = 8'h00;
reg_space[1112] = 8'h00;
reg_space[1113] = 8'h00;
reg_space[1114] = 8'h00;
reg_space[1115] = 8'h00;
reg_space[1116] = 8'h00;
reg_space[1117] = 8'h00;
reg_space[1118] = 8'h00;
reg_space[1119] = 8'h00;
reg_space[1120] = 8'h00;
reg_space[1121] = 8'h00;
reg_space[1122] = 8'h00;
reg_space[1123] = 8'h00;
reg_space[1124] = 8'h00;
reg_space[1125] = 8'h00;
reg_space[1126] = 8'h00;
reg_space[1127] = 8'h00;
reg_space[1128] = 8'h00;
reg_space[1129] = 8'h00;
reg_space[1130] = 8'h00;
reg_space[1131] = 8'h00;
reg_space[1132] = 8'h00;
reg_space[1133] = 8'h00;
reg_space[1134] = 8'h00;
reg_space[1135] = 8'h00;
reg_space[1136] = 8'h00;
reg_space[1137] = 8'h00;
reg_space[1138] = 8'h00;
reg_space[1139] = 8'h00;
reg_space[1140] = 8'h00;
reg_space[1141] = 8'h00;
reg_space[1142] = 8'h00;
reg_space[1143] = 8'h00;
reg_space[1144] = 8'h00;
reg_space[1145] = 8'h00;
reg_space[1146] = 8'h00;
reg_space[1147] = 8'h00;
reg_space[1148] = 8'h00;
reg_space[1149] = 8'h00;
reg_space[1150] = 8'h00;
reg_space[1151] = 8'h00;
reg_space[1152] = 8'h00;
reg_space[1153] = 8'h00;
reg_space[1154] = 8'h00;
reg_space[1155] = 8'h00;
reg_space[1156] = 8'h00;
reg_space[1157] = 8'h00;
reg_space[1158] = 8'h00;
reg_space[1159] = 8'h00;
reg_space[1160] = 8'h00;
reg_space[1161] = 8'h00;
reg_space[1162] = 8'h00;
reg_space[1163] = 8'h00;
reg_space[1164] = 8'h00;
reg_space[1165] = 8'h00;
reg_space[1166] = 8'h00;
reg_space[1167] = 8'h00;
reg_space[1168] = 8'h00;
reg_space[1169] = 8'h00;
reg_space[1170] = 8'h00;
reg_space[1171] = 8'h00;
reg_space[1172] = 8'h00;
reg_space[1173] = 8'h00;
reg_space[1174] = 8'h00;
reg_space[1175] = 8'h00;
reg_space[1176] = 8'h00;
reg_space[1177] = 8'h00;
reg_space[1178] = 8'h00;
reg_space[1179] = 8'h00;
reg_space[1180] = 8'h00;
reg_space[1181] = 8'h00;
reg_space[1182] = 8'h00;
reg_space[1183] = 8'h00;
reg_space[1184] = 8'h00;
reg_space[1185] = 8'h00;
reg_space[1186] = 8'h00;
reg_space[1187] = 8'h00;
reg_space[1188] = 8'h00;
reg_space[1189] = 8'h00;
reg_space[1190] = 8'h00;
reg_space[1191] = 8'h00;
reg_space[1192] = 8'h00;
reg_space[1193] = 8'h00;
reg_space[1194] = 8'h00;
reg_space[1195] = 8'h00;
reg_space[1196] = 8'h00;
reg_space[1197] = 8'h00;
reg_space[1198] = 8'h00;
reg_space[1199] = 8'h00;
reg_space[1200] = 8'h00;
reg_space[1201] = 8'h00;
reg_space[1202] = 8'h00;
reg_space[1203] = 8'h00;
reg_space[1204] = 8'h00;
reg_space[1205] = 8'h00;
reg_space[1206] = 8'h00;
reg_space[1207] = 8'h00;
reg_space[1208] = 8'h00;
reg_space[1209] = 8'h00;
reg_space[1210] = 8'h00;
reg_space[1211] = 8'h00;
reg_space[1212] = 8'h00;
reg_space[1213] = 8'h00;
reg_space[1214] = 8'h00;
reg_space[1215] = 8'h00;
reg_space[1216] = 8'h00;
reg_space[1217] = 8'h00;
reg_space[1218] = 8'h00;
reg_space[1219] = 8'h00;
reg_space[1220] = 8'h00;
reg_space[1221] = 8'h00;
reg_space[1222] = 8'h00;
reg_space[1223] = 8'h00;
reg_space[1224] = 8'h00;
reg_space[1225] = 8'h00;
reg_space[1226] = 8'h00;
reg_space[1227] = 8'h00;
reg_space[1228] = 8'h00;
reg_space[1229] = 8'h00;
reg_space[1230] = 8'h00;
reg_space[1231] = 8'h00;
reg_space[1232] = 8'h00;
reg_space[1233] = 8'h00;
reg_space[1234] = 8'h00;
reg_space[1235] = 8'h00;
reg_space[1236] = 8'h00;
reg_space[1237] = 8'h00;
reg_space[1238] = 8'h00;
reg_space[1239] = 8'h00;
reg_space[1240] = 8'h00;
reg_space[1241] = 8'h00;
reg_space[1242] = 8'h00;
reg_space[1243] = 8'h00;
reg_space[1244] = 8'h00;
reg_space[1245] = 8'h00;
reg_space[1246] = 8'h00;
reg_space[1247] = 8'h00;
reg_space[1248] = 8'h00;
reg_space[1249] = 8'h00;
reg_space[1250] = 8'h00;
reg_space[1251] = 8'h00;
reg_space[1252] = 8'h00;
reg_space[1253] = 8'h00;
reg_space[1254] = 8'h00;
reg_space[1255] = 8'h00;
reg_space[1256] = 8'h00;
reg_space[1257] = 8'h00;
reg_space[1258] = 8'h00;
reg_space[1259] = 8'h00;
reg_space[1260] = 8'h00;
reg_space[1261] = 8'h00;
reg_space[1262] = 8'h00;
reg_space[1263] = 8'h00;
reg_space[1264] = 8'h00;
reg_space[1265] = 8'h00;
reg_space[1266] = 8'h00;
reg_space[1267] = 8'h00;
reg_space[1268] = 8'h00;
reg_space[1269] = 8'h00;
reg_space[1270] = 8'h00;
reg_space[1271] = 8'h00;
reg_space[1272] = 8'h00;
reg_space[1273] = 8'h00;
reg_space[1274] = 8'h00;
reg_space[1275] = 8'h00;
reg_space[1276] = 8'h00;
reg_space[1277] = 8'h00;
reg_space[1278] = 8'h00;
reg_space[1279] = 8'h00;
reg_space[1280] = 8'h00;
reg_space[1281] = 8'h00;
reg_space[1282] = 8'h00;
reg_space[1283] = 8'h00;
reg_space[1284] = 8'h00;
reg_space[1285] = 8'h00;
reg_space[1286] = 8'h00;
reg_space[1287] = 8'h00;
reg_space[1288] = 8'h00;
reg_space[1289] = 8'h00;
reg_space[1290] = 8'h00;
reg_space[1291] = 8'h00;
reg_space[1292] = 8'h00;
reg_space[1293] = 8'h00;
reg_space[1294] = 8'h00;
reg_space[1295] = 8'h00;
reg_space[1296] = 8'h00;
reg_space[1297] = 8'h00;
reg_space[1298] = 8'h00;
reg_space[1299] = 8'h00;
reg_space[1300] = 8'h00;
reg_space[1301] = 8'h00;
reg_space[1302] = 8'h00;
reg_space[1303] = 8'h00;
reg_space[1304] = 8'h00;
reg_space[1305] = 8'h00;
reg_space[1306] = 8'h00;
reg_space[1307] = 8'h00;
reg_space[1308] = 8'h00;
reg_space[1309] = 8'h00;
reg_space[1310] = 8'h00;
reg_space[1311] = 8'h00;
reg_space[1312] = 8'h00;
reg_space[1313] = 8'h00;
reg_space[1314] = 8'h00;
reg_space[1315] = 8'h00;
reg_space[1316] = 8'h00;
reg_space[1317] = 8'h00;
reg_space[1318] = 8'h00;
reg_space[1319] = 8'h00;
reg_space[1320] = 8'h00;
reg_space[1321] = 8'h00;
reg_space[1322] = 8'h00;
reg_space[1323] = 8'h00;
reg_space[1324] = 8'h00;
reg_space[1325] = 8'h00;
reg_space[1326] = 8'h00;
reg_space[1327] = 8'h00;
reg_space[1328] = 8'h00;
reg_space[1329] = 8'h00;
reg_space[1330] = 8'h00;
reg_space[1331] = 8'h00;
reg_space[1332] = 8'h00;
reg_space[1333] = 8'h00;
reg_space[1334] = 8'h00;
reg_space[1335] = 8'h00;
reg_space[1336] = 8'h00;
reg_space[1337] = 8'h00;
reg_space[1338] = 8'h00;
reg_space[1339] = 8'h00;
reg_space[1340] = 8'h00;
reg_space[1341] = 8'h00;
reg_space[1342] = 8'h00;
reg_space[1343] = 8'h00;
reg_space[1344] = 8'h00;
reg_space[1345] = 8'h00;
reg_space[1346] = 8'h00;
reg_space[1347] = 8'h00;
reg_space[1348] = 8'h00;
reg_space[1349] = 8'h00;
reg_space[1350] = 8'h00;
reg_space[1351] = 8'h00;
reg_space[1352] = 8'h00;
reg_space[1353] = 8'h00;
reg_space[1354] = 8'h00;
reg_space[1355] = 8'h00;
reg_space[1356] = 8'h00;
reg_space[1357] = 8'h00;
reg_space[1358] = 8'h00;
reg_space[1359] = 8'h00;
reg_space[1360] = 8'h00;
reg_space[1361] = 8'h00;
reg_space[1362] = 8'h00;
reg_space[1363] = 8'h00;
reg_space[1364] = 8'h00;
reg_space[1365] = 8'h00;
reg_space[1366] = 8'h00;
reg_space[1367] = 8'h00;
reg_space[1368] = 8'h00;
reg_space[1369] = 8'h00;
reg_space[1370] = 8'h00;
reg_space[1371] = 8'h00;
reg_space[1372] = 8'h00;
reg_space[1373] = 8'h00;
reg_space[1374] = 8'h00;
reg_space[1375] = 8'h00;
reg_space[1376] = 8'h00;
reg_space[1377] = 8'h00;
reg_space[1378] = 8'h00;
reg_space[1379] = 8'h00;
reg_space[1380] = 8'h00;
reg_space[1381] = 8'h00;
reg_space[1382] = 8'h00;
reg_space[1383] = 8'h00;
reg_space[1384] = 8'h00;
reg_space[1385] = 8'h00;
reg_space[1386] = 8'h00;
reg_space[1387] = 8'h00;
reg_space[1388] = 8'h00;
reg_space[1389] = 8'h00;
reg_space[1390] = 8'h00;
reg_space[1391] = 8'h00;
reg_space[1392] = 8'h00;
reg_space[1393] = 8'h00;
reg_space[1394] = 8'h00;
reg_space[1395] = 8'h00;
reg_space[1396] = 8'h00;
reg_space[1397] = 8'h00;
reg_space[1398] = 8'h00;
reg_space[1399] = 8'h00;
reg_space[1400] = 8'h00;
reg_space[1401] = 8'h00;
reg_space[1402] = 8'h00;
reg_space[1403] = 8'h00;
reg_space[1404] = 8'h00;
reg_space[1405] = 8'h00;
reg_space[1406] = 8'h00;
reg_space[1407] = 8'h00;
reg_space[1408] = 8'h00;
reg_space[1409] = 8'h00;
reg_space[1410] = 8'h00;
reg_space[1411] = 8'h00;
reg_space[1412] = 8'h00;
reg_space[1413] = 8'h00;
reg_space[1414] = 8'h00;
reg_space[1415] = 8'h00;
reg_space[1416] = 8'h00;
reg_space[1417] = 8'h00;
reg_space[1418] = 8'h00;
reg_space[1419] = 8'h00;
reg_space[1420] = 8'h00;
reg_space[1421] = 8'h00;
reg_space[1422] = 8'h00;
reg_space[1423] = 8'h00;
reg_space[1424] = 8'h00;
reg_space[1425] = 8'h00;
reg_space[1426] = 8'h00;
reg_space[1427] = 8'h00;
reg_space[1428] = 8'h00;
reg_space[1429] = 8'h00;
reg_space[1430] = 8'h00;
reg_space[1431] = 8'h00;
reg_space[1432] = 8'h00;
reg_space[1433] = 8'h00;
reg_space[1434] = 8'h00;
reg_space[1435] = 8'h00;
reg_space[1436] = 8'h00;
reg_space[1437] = 8'h00;
reg_space[1438] = 8'h00;
reg_space[1439] = 8'h00;
reg_space[1440] = 8'h00;
reg_space[1441] = 8'h00;
reg_space[1442] = 8'h00;
reg_space[1443] = 8'h00;
reg_space[1444] = 8'h00;
reg_space[1445] = 8'h00;
reg_space[1446] = 8'h00;
reg_space[1447] = 8'h00;
reg_space[1448] = 8'h00;
reg_space[1449] = 8'h00;
reg_space[1450] = 8'h00;
reg_space[1451] = 8'h00;
reg_space[1452] = 8'h00;
reg_space[1453] = 8'h00;
reg_space[1454] = 8'h00;
reg_space[1455] = 8'h00;
reg_space[1456] = 8'h00;
reg_space[1457] = 8'h00;
reg_space[1458] = 8'h00;
reg_space[1459] = 8'h00;
reg_space[1460] = 8'h00;
reg_space[1461] = 8'h00;
reg_space[1462] = 8'h00;
reg_space[1463] = 8'h00;
reg_space[1464] = 8'h00;
reg_space[1465] = 8'h00;
reg_space[1466] = 8'h00;
reg_space[1467] = 8'h00;
reg_space[1468] = 8'h00;
reg_space[1469] = 8'h00;
reg_space[1470] = 8'h00;
reg_space[1471] = 8'h00;
reg_space[1472] = 8'h00;
reg_space[1473] = 8'h00;
reg_space[1474] = 8'h00;
reg_space[1475] = 8'h00;
reg_space[1476] = 8'h00;
reg_space[1477] = 8'h00;
reg_space[1478] = 8'h00;
reg_space[1479] = 8'h00;
reg_space[1480] = 8'h00;
reg_space[1481] = 8'h00;
reg_space[1482] = 8'h00;
reg_space[1483] = 8'h00;
reg_space[1484] = 8'h00;
reg_space[1485] = 8'h00;
reg_space[1486] = 8'h00;
reg_space[1487] = 8'h00;
reg_space[1488] = 8'h00;
reg_space[1489] = 8'h00;
reg_space[1490] = 8'h00;
reg_space[1491] = 8'h00;
reg_space[1492] = 8'h00;
reg_space[1493] = 8'h00;
reg_space[1494] = 8'h00;
reg_space[1495] = 8'h00;
reg_space[1496] = 8'h00;
reg_space[1497] = 8'h00;
reg_space[1498] = 8'h00;
reg_space[1499] = 8'h00;
reg_space[1500] = 8'h00;
reg_space[1501] = 8'h00;
reg_space[1502] = 8'h00;
reg_space[1503] = 8'h00;
reg_space[1504] = 8'h00;
reg_space[1505] = 8'h00;
reg_space[1506] = 8'h00;
reg_space[1507] = 8'h00;
reg_space[1508] = 8'h00;
reg_space[1509] = 8'h00;
reg_space[1510] = 8'h00;
reg_space[1511] = 8'h00;
reg_space[1512] = 8'h00;
reg_space[1513] = 8'h00;
reg_space[1514] = 8'h00;
reg_space[1515] = 8'h00;
reg_space[1516] = 8'h00;
reg_space[1517] = 8'h00;
reg_space[1518] = 8'h00;
reg_space[1519] = 8'h00;
reg_space[1520] = 8'h00;
reg_space[1521] = 8'h00;
reg_space[1522] = 8'h00;
reg_space[1523] = 8'h00;
reg_space[1524] = 8'h00;
reg_space[1525] = 8'h00;
reg_space[1526] = 8'h00;
reg_space[1527] = 8'h00;
reg_space[1528] = 8'h00;
reg_space[1529] = 8'h00;
reg_space[1530] = 8'h00;
reg_space[1531] = 8'h00;
reg_space[1532] = 8'h00;
reg_space[1533] = 8'h00;
reg_space[1534] = 8'h00;
reg_space[1535] = 8'h00;
reg_space[1536] = 8'h00;
reg_space[1537] = 8'h00;
reg_space[1538] = 8'h00;
reg_space[1539] = 8'h00;
reg_space[1540] = 8'h00;
reg_space[1541] = 8'h00;
reg_space[1542] = 8'h00;
reg_space[1543] = 8'h00;
reg_space[1544] = 8'h00;
reg_space[1545] = 8'h00;
reg_space[1546] = 8'h00;
reg_space[1547] = 8'h00;
reg_space[1548] = 8'h00;
reg_space[1549] = 8'h00;
reg_space[1550] = 8'h00;
reg_space[1551] = 8'h00;
reg_space[1552] = 8'h00;
reg_space[1553] = 8'h00;
reg_space[1554] = 8'h00;
reg_space[1555] = 8'h00;
reg_space[1556] = 8'h00;
reg_space[1557] = 8'h00;
reg_space[1558] = 8'h00;
reg_space[1559] = 8'h00;
reg_space[1560] = 8'h00;
reg_space[1561] = 8'h00;
reg_space[1562] = 8'h00;
reg_space[1563] = 8'h00;
reg_space[1564] = 8'h00;
reg_space[1565] = 8'h00;
reg_space[1566] = 8'h00;
reg_space[1567] = 8'h00;
reg_space[1568] = 8'h00;
reg_space[1569] = 8'h00;
reg_space[1570] = 8'h00;
reg_space[1571] = 8'h00;
reg_space[1572] = 8'h00;
reg_space[1573] = 8'h00;
reg_space[1574] = 8'h00;
reg_space[1575] = 8'h00;
reg_space[1576] = 8'h00;
reg_space[1577] = 8'h00;
reg_space[1578] = 8'h00;
reg_space[1579] = 8'h00;
reg_space[1580] = 8'h00;
reg_space[1581] = 8'h00;
reg_space[1582] = 8'h00;
reg_space[1583] = 8'h00;
reg_space[1584] = 8'h00;
reg_space[1585] = 8'h00;
reg_space[1586] = 8'h00;
reg_space[1587] = 8'h00;
reg_space[1588] = 8'h00;
reg_space[1589] = 8'h00;
reg_space[1590] = 8'h00;
reg_space[1591] = 8'h00;
reg_space[1592] = 8'h00;
reg_space[1593] = 8'h00;
reg_space[1594] = 8'h00;
reg_space[1595] = 8'h00;
reg_space[1596] = 8'h00;
reg_space[1597] = 8'h00;
reg_space[1598] = 8'h00;
reg_space[1599] = 8'h00;
reg_space[1600; = 8'h00;
reg_space[1601] = 8'h00;
reg_space[1602] = 8'h00;
reg_space[1603] = 8'h00;
reg_space[1604] = 8'h00;
reg_space[1605] = 8'h00;
reg_space[1606] = 8'h00;
reg_space[1607] = 8'h00;
reg_space[1608] = 8'h00;
reg_space[1609] = 8'h00;
reg_space[1610] = 8'h00;
reg_space[1611] = 8'h00;
reg_space[1612] = 8'h00;
reg_space[1613] = 8'h00;
reg_space[1614] = 8'h00;
reg_space[1615] = 8'h00;
reg_space[1616] = 8'h00;
reg_space[1617] = 8'h00;
reg_space[1618] = 8'h00;
reg_space[1619] = 8'h00;
reg_space[1620] = 8'h00;
reg_space[1621] = 8'h00;
reg_space[1622] = 8'h00;
reg_space[1623] = 8'h00;
reg_space[1624] = 8'h00;
reg_space[1625] = 8'h00;
reg_space[1626] = 8'h00;
reg_space[1627] = 8'h00;
reg_space[1628] = 8'h00;
reg_space[1629] = 8'h00;
reg_space[1630] = 8'h00;
reg_space[1631] = 8'h00;
reg_space[1632] = 8'h00;
reg_space[1633] = 8'h00;
reg_space[1634] = 8'h00;
reg_space[1635] = 8'h00;
reg_space[1636] = 8'h00;
reg_space[1637] = 8'h00;
reg_space[1638] = 8'h00;
reg_space[1639] = 8'h00;
reg_space[1640] = 8'h00;
reg_space[1641] = 8'h00;
reg_space[1642] = 8'h00;
reg_space[1643] = 8'h00;
reg_space[1644] = 8'h00;
reg_space[1645] = 8'h00;
reg_space[1646] = 8'h00;
reg_space[1647] = 8'h00;
reg_space[1648] = 8'h00;
reg_space[1649] = 8'h00;
reg_space[1650] = 8'h00;
reg_space[1651] = 8'h00;
reg_space[1652] = 8'h00;
reg_space[1653] = 8'h00;
reg_space[1654] = 8'h00;
reg_space[1655] = 8'h00;
reg_space[1656] = 8'h00;
reg_space[1657] = 8'h00;
reg_space[1658] = 8'h00;
reg_space[1659] = 8'h00;
reg_space[1660] = 8'h00;
reg_space[1661] = 8'h00;
reg_space[1662] = 8'h00;
reg_space[1663] = 8'h00;
reg_space[1664] = 8'h00;
reg_space[1665] = 8'h00;
reg_space[1666] = 8'h00;
reg_space[1667] = 8'h00;
reg_space[1668] = 8'h00;
reg_space[1669] = 8'h00;
reg_space[1670] = 8'h00;
reg_space[1671] = 8'h00;
reg_space[1672] = 8'h00;
reg_space[1673] = 8'h00;
reg_space[1674] = 8'h00;
reg_space[1675] = 8'h00;
reg_space[1676] = 8'h00;
reg_space[1677] = 8'h00;
reg_space[1678] = 8'h00;
reg_space[1679] = 8'h00;
reg_space[1680] = 8'h00;
reg_space[1681] = 8'h00;
reg_space[1682] = 8'h00;
reg_space[1683] = 8'h00;
reg_space[1684] = 8'h00;
reg_space[1685] = 8'h00;
reg_space[1686] = 8'h00;
reg_space[1687] = 8'h00;
reg_space[1688] = 8'h00;
reg_space[1689] = 8'h00;
reg_space[1690] = 8'h00;
reg_space[1691] = 8'h00;
reg_space[1692] = 8'h00;
reg_space[1693] = 8'h00;
reg_space[1694] = 8'h00;
reg_space[1695] = 8'h00;
reg_space[1696] = 8'h00;
reg_space[1697] = 8'h00;
reg_space[1698] = 8'h00;
reg_space[1699] = 8'h00;
reg_space[1700; = 8'h00;
reg_space[1701] = 8'h00;
reg_space[1702] = 8'h00;
reg_space[1703] = 8'h00;
reg_space[1704] = 8'h00;
reg_space[1705] = 8'h00;
reg_space[1706] = 8'h00;
reg_space[1707] = 8'h00;
reg_space[1708] = 8'h00;
reg_space[1709] = 8'h00;
reg_space[1710] = 8'h00;
reg_space[1711] = 8'h00;
reg_space[1712] = 8'h00;
reg_space[1713] = 8'h00;
reg_space[1714] = 8'h00;
reg_space[1715] = 8'h00;
reg_space[1716] = 8'h00;
reg_space[1717] = 8'h00;
reg_space[1718] = 8'h00;
reg_space[1719] = 8'h00;
reg_space[1720] = 8'h00;
reg_space[1721] = 8'h00;
reg_space[1722] = 8'h00;
reg_space[1723] = 8'h00;
reg_space[1724] = 8'h00;
reg_space[1725] = 8'h00;
reg_space[1726] = 8'h00;
reg_space[1727] = 8'h00;
reg_space[1728] = 8'h00;
reg_space[1729] = 8'h00;
reg_space[1730] = 8'h00;
reg_space[1731] = 8'h00;
reg_space[1732] = 8'h00;
reg_space[1733] = 8'h00;
reg_space[1734] = 8'h00;
reg_space[1735] = 8'h00;
reg_space[1736] = 8'h00;
reg_space[1737] = 8'h00;
reg_space[1738] = 8'h00;
reg_space[1739] = 8'h00;
reg_space[1740] = 8'h00;
reg_space[1741] = 8'h00;
reg_space[1742] = 8'h00;
reg_space[1743] = 8'h00;
reg_space[1744] = 8'h00;
reg_space[1745] = 8'h00;
reg_space[1746] = 8'h00;
reg_space[1747] = 8'h00;
reg_space[1748] = 8'h00;
reg_space[1749] = 8'h00;
reg_space[1750] = 8'h00;
reg_space[1751] = 8'h00;
reg_space[1752] = 8'h00;
reg_space[1753] = 8'h00;
reg_space[1754] = 8'h00;
reg_space[1755] = 8'h00;
reg_space[1756] = 8'h00;
reg_space[1757] = 8'h00;
reg_space[1758] = 8'h00;
reg_space[1759] = 8'h00;
reg_space[1760] = 8'h00;
reg_space[1761] = 8'h00;
reg_space[1762] = 8'h00;
reg_space[1763] = 8'h00;
reg_space[1764] = 8'h00;
reg_space[1765] = 8'h00;
reg_space[1766] = 8'h00;
reg_space[1767] = 8'h00;
reg_space[1768] = 8'h00;
reg_space[1769] = 8'h00;
reg_space[1770] = 8'h00;
reg_space[1771] = 8'h00;
reg_space[1772] = 8'h00;
reg_space[1773] = 8'h00;
reg_space[1774] = 8'h00;
reg_space[1775] = 8'h00;
reg_space[1776] = 8'h00;
reg_space[1777] = 8'h00;
reg_space[1778] = 8'h00;
reg_space[1779] = 8'h00;
reg_space[1780] = 8'h00;
reg_space[1781] = 8'h00;
reg_space[1782] = 8'h00;
reg_space[1783] = 8'h00;
reg_space[1784] = 8'h00;
reg_space[1785] = 8'h00;
reg_space[1786] = 8'h00;
reg_space[1787] = 8'h00;
reg_space[1788] = 8'h00;
reg_space[1789] = 8'h00;
reg_space[1790] = 8'h00;
reg_space[1791] = 8'h00;
reg_space[1792] = 8'h00;
reg_space[1793] = 8'h00;
reg_space[1794] = 8'h00;
reg_space[1795] = 8'h00;
reg_space[1796] = 8'h00;
reg_space[1797] = 8'h00;
reg_space[1798] = 8'h00;
reg_space[1799] = 8'h00;
reg_space[1800; = 8'h00;
reg_space[1801] = 8'h00;
reg_space[1802] = 8'h00;
reg_space[1803] = 8'h00;
reg_space[1804] = 8'h00;
reg_space[1805] = 8'h00;
reg_space[1806] = 8'h00;
reg_space[1807] = 8'h00;
reg_space[1808] = 8'h00;
reg_space[1809] = 8'h00;
reg_space[1810] = 8'h00;
reg_space[1811] = 8'h00;
reg_space[1812] = 8'h00;
reg_space[1813] = 8'h00;
reg_space[1814] = 8'h00;
reg_space[1815] = 8'h00;
reg_space[1816] = 8'h00;
reg_space[1817] = 8'h00;
reg_space[1818] = 8'h00;
reg_space[1819] = 8'h00;
reg_space[1820] = 8'h00;
reg_space[1821] = 8'h00;
reg_space[1822] = 8'h00;
reg_space[1823] = 8'h00;
reg_space[1824] = 8'h00;
reg_space[1825] = 8'h00;
reg_space[1826] = 8'h00;
reg_space[1827] = 8'h00;
reg_space[1828] = 8'h00;
reg_space[1829] = 8'h00;
reg_space[1830] = 8'h00;
reg_space[1831] = 8'h00;
reg_space[1832] = 8'h00;
reg_space[1833] = 8'h00;
reg_space[1834] = 8'h00;
reg_space[1835] = 8'h00;
reg_space[1836] = 8'h00;
reg_space[1837] = 8'h00;
reg_space[1838] = 8'h00;
reg_space[1839] = 8'h00;
reg_space[1840] = 8'h00;
reg_space[1841] = 8'h00;
reg_space[1842] = 8'h00;
reg_space[1843] = 8'h00;
reg_space[1844] = 8'h00;
reg_space[1845] = 8'h00;
reg_space[1846] = 8'h00;
reg_space[1847] = 8'h00;
reg_space[1848] = 8'h00;
reg_space[1849] = 8'h00;
reg_space[1850] = 8'h00;
reg_space[1851] = 8'h00;
reg_space[1852] = 8'h00;
reg_space[1853] = 8'h00;
reg_space[1854] = 8'h00;
reg_space[1855] = 8'h00;
reg_space[1856] = 8'h00;
reg_space[1857] = 8'h00;
reg_space[1858] = 8'h00;
reg_space[1859] = 8'h00;
reg_space[1860] = 8'h00;
reg_space[1861] = 8'h00;
reg_space[1862] = 8'h00;
reg_space[1863] = 8'h00;
reg_space[1864] = 8'h00;
reg_space[1865] = 8'h00;
reg_space[1866] = 8'h00;
reg_space[1867] = 8'h00;
reg_space[1868] = 8'h00;
reg_space[1869] = 8'h00;
reg_space[1870] = 8'h00;
reg_space[1871] = 8'h00;
reg_space[1872] = 8'h00;
reg_space[1873] = 8'h00;
reg_space[1874] = 8'h00;
reg_space[1875] = 8'h00;
reg_space[1876] = 8'h00;
reg_space[1877] = 8'h00;
reg_space[1878] = 8'h00;
reg_space[1879] = 8'h00;
reg_space[1880] = 8'h00;
reg_space[1881] = 8'h00;
reg_space[1882] = 8'h00;
reg_space[1883] = 8'h00;
reg_space[1884] = 8'h00;
reg_space[1885] = 8'h00;
reg_space[1886] = 8'h00;
reg_space[1887] = 8'h00;
reg_space[1888] = 8'h00;
reg_space[1889] = 8'h00;
reg_space[1890] = 8'h00;
reg_space[1891] = 8'h00;
reg_space[1892] = 8'h00;
reg_space[1893] = 8'h00;
reg_space[1894] = 8'h00;
reg_space[1895] = 8'h00;
reg_space[1896] = 8'h00;
reg_space[1897] = 8'h00;
reg_space[1898] = 8'h00;
reg_space[1899] = 8'h00;
reg_space[1900; = 8'h00;
reg_space[1901] = 8'h00;
reg_space[1902] = 8'h00;
reg_space[1903] = 8'h00;
reg_space[1904] = 8'h00;
reg_space[1905] = 8'h00;
reg_space[1906] = 8'h00;
reg_space[1907] = 8'h00;
reg_space[1908] = 8'h00;
reg_space[1909] = 8'h00;
reg_space[1910] = 8'h00;
reg_space[1911] = 8'h00;
reg_space[1912] = 8'h00;
reg_space[1913] = 8'h00;
reg_space[1914] = 8'h00;
reg_space[1915] = 8'h00;
reg_space[1916] = 8'h00;
reg_space[1917] = 8'h00;
reg_space[1918] = 8'h00;
reg_space[1919] = 8'h00;
reg_space[1920] = 8'h00;
reg_space[1921] = 8'h00;
reg_space[1922] = 8'h00;
reg_space[1923] = 8'h00;
reg_space[1924] = 8'h00;
reg_space[1925] = 8'h00;
reg_space[1926] = 8'h00;
reg_space[1927] = 8'h00;
reg_space[1928] = 8'h00;
reg_space[1929] = 8'h00;
reg_space[1930] = 8'h00;
reg_space[1931] = 8'h00;
reg_space[1932] = 8'h00;
reg_space[1933] = 8'h00;
reg_space[1934] = 8'h00;
reg_space[1935] = 8'h00;
reg_space[1936] = 8'h00;
reg_space[1937] = 8'h00;
reg_space[1938] = 8'h00;
reg_space[1939] = 8'h00;
reg_space[1940] = 8'h00;
reg_space[1941] = 8'h00;
reg_space[1942] = 8'h00;
reg_space[1943] = 8'h00;
reg_space[1944] = 8'h00;
reg_space[1945] = 8'h00;
reg_space[1946] = 8'h00;
reg_space[1947] = 8'h00;
reg_space[1948] = 8'h00;
reg_space[1949] = 8'h00;
reg_space[1950] = 8'h00;
reg_space[1951] = 8'h00;
reg_space[1952] = 8'h00;
reg_space[1953] = 8'h00;
reg_space[1954] = 8'h00;
reg_space[1955] = 8'h00;
reg_space[1956] = 8'h00;
reg_space[1957] = 8'h00;
reg_space[1958] = 8'h00;
reg_space[1959] = 8'h00;
reg_space[1960] = 8'h00;
reg_space[1961] = 8'h00;
reg_space[1962] = 8'h00;
reg_space[1963] = 8'h00;
reg_space[1964] = 8'h00;
reg_space[1965] = 8'h00;
reg_space[1966] = 8'h00;
reg_space[1967] = 8'h00;
reg_space[1968] = 8'h00;
reg_space[1969] = 8'h00;
reg_space[1970] = 8'h00;
reg_space[1971] = 8'h00;
reg_space[1972] = 8'h00;
reg_space[1973] = 8'h00;
reg_space[1974] = 8'h00;
reg_space[1975] = 8'h00;
reg_space[1976] = 8'h00;
reg_space[1977] = 8'h00;
reg_space[1978] = 8'h00;
reg_space[1979] = 8'h00;
reg_space[1980] = 8'h00;
reg_space[1981] = 8'h00;
reg_space[1982] = 8'h00;
reg_space[1983] = 8'h00;
reg_space[1984] = 8'h00;
reg_space[1985] = 8'h00;
reg_space[1986] = 8'h00;
reg_space[1987] = 8'h00;
reg_space[1988] = 8'h00;
reg_space[1989] = 8'h00;
reg_space[1990] = 8'h00;
reg_space[1991] = 8'h00;
reg_space[1992] = 8'h00;
reg_space[1993] = 8'h00;
reg_space[1994] = 8'h00;
reg_space[1995] = 8'h00;
reg_space[1996] = 8'h00;
reg_space[1997] = 8'h00;
reg_space[1998] = 8'h00;
reg_space[1999] = 8'h00;
reg_space[200;0] = 8'h00;
reg_space[200;1] = 8'h00;
reg_space[200;2] = 8'h00;
reg_space[200;3] = 8'h00;
reg_space[200;4] = 8'h00;
reg_space[200;5] = 8'h00;
reg_space[200;6] = 8'h00;
reg_space[200;7] = 8'h00;
reg_space[200;8] = 8'h00;
reg_space[200;9] = 8'h00;
reg_space[2010] = 8'h00;
reg_space[2011] = 8'h00;
reg_space[2012] = 8'h00;
reg_space[2013] = 8'h00;
reg_space[2014] = 8'h00;
reg_space[2015] = 8'h00;
reg_space[2016] = 8'h00;
reg_space[2017] = 8'h00;
reg_space[2018] = 8'h00;
reg_space[2019] = 8'h00;
reg_space[2020] = 8'h00;
reg_space[2021] = 8'h00;
reg_space[2022] = 8'h00;
reg_space[2023] = 8'h00;
reg_space[2024] = 8'h00;
reg_space[2025] = 8'h00;
reg_space[2026] = 8'h00;
reg_space[2027] = 8'h00;
reg_space[2028] = 8'h00;
reg_space[2029] = 8'h00;
reg_space[2030] = 8'h00;
reg_space[2031] = 8'h00;
reg_space[2032] = 8'h00;
reg_space[2033] = 8'h00;
reg_space[2034] = 8'h00;
reg_space[2035] = 8'h00;
reg_space[2036] = 8'h00;
reg_space[2037] = 8'h00;
reg_space[2038] = 8'h00;
reg_space[2039] = 8'h00;
reg_space[2040] = 8'h00;
reg_space[2041] = 8'h00;
reg_space[2042] = 8'h00;
reg_space[2043] = 8'h00;
reg_space[2044] = 8'h00;
reg_space[2045] = 8'h00;
reg_space[2046] = 8'h00;
reg_space[2047] = 8'h00;
reg_space[2048] = 8'h00;
reg_space[2049] = 8'h00;
reg_space[2050] = 8'h00;
reg_space[2051] = 8'h00;
reg_space[2052] = 8'h00;
reg_space[2053] = 8'h00;
reg_space[2054] = 8'h00;
reg_space[2055] = 8'h00;
reg_space[2056] = 8'h00;
reg_space[2057] = 8'h00;
reg_space[2058] = 8'h00;
reg_space[2059] = 8'h00;
reg_space[2060] = 8'h00;
reg_space[2061] = 8'h00;
reg_space[2062] = 8'h00;
reg_space[2063] = 8'h00;
reg_space[2064] = 8'h00;
reg_space[2065] = 8'h00;
reg_space[2066] = 8'h00;
reg_space[2067] = 8'h00;
reg_space[2068] = 8'h00;
reg_space[2069] = 8'h00;
reg_space[2070] = 8'h00;
reg_space[2071] = 8'h00;
reg_space[2072] = 8'h00;
reg_space[2073] = 8'h00;
reg_space[2074] = 8'h00;
reg_space[2075] = 8'h00;
reg_space[2076] = 8'h00;
reg_space[2077] = 8'h00;
reg_space[2078] = 8'h00;
reg_space[2079] = 8'h00;
reg_space[2080] = 8'h00;
reg_space[2081] = 8'h00;
reg_space[2082] = 8'h00;
reg_space[2083] = 8'h00;
reg_space[2084] = 8'h00;
reg_space[2085] = 8'h00;
reg_space[2086] = 8'h00;
reg_space[2087] = 8'h00;
reg_space[2088] = 8'h00;
reg_space[2089] = 8'h00;
reg_space[2090] = 8'h00;
reg_space[2091] = 8'h00;
reg_space[2092] = 8'h00;
reg_space[2093] = 8'h00;
reg_space[2094] = 8'h00;
reg_space[2095] = 8'h00;
reg_space[2096] = 8'h00;
reg_space[2097] = 8'h00;
reg_space[2098] = 8'h00;
reg_space[2099] = 8'h00;
reg_space[2100; = 8'h00;
reg_space[2101] = 8'h00;
reg_space[2102] = 8'h00;
reg_space[2103] = 8'h00;
reg_space[2104] = 8'h00;
reg_space[2105] = 8'h00;
reg_space[2106] = 8'h00;
reg_space[2107] = 8'h00;
reg_space[2108] = 8'h00;
reg_space[2109] = 8'h00;
reg_space[2110] = 8'h00;
reg_space[2111] = 8'h00;
reg_space[2112] = 8'h00;
reg_space[2113] = 8'h00;
reg_space[2114] = 8'h00;
reg_space[2115] = 8'h00;
reg_space[2116] = 8'h00;
reg_space[2117] = 8'h00;
reg_space[2118] = 8'h00;
reg_space[2119] = 8'h00;
reg_space[2120] = 8'h00;
reg_space[2121] = 8'h00;
reg_space[2122] = 8'h00;
reg_space[2123] = 8'h00;
reg_space[2124] = 8'h00;
reg_space[2125] = 8'h00;
reg_space[2126] = 8'h00;
reg_space[2127] = 8'h00;
reg_space[2128] = 8'h00;
reg_space[2129] = 8'h00;
reg_space[2130] = 8'h00;
reg_space[2131] = 8'h00;
reg_space[2132] = 8'h00;
reg_space[2133] = 8'h00;
reg_space[2134] = 8'h00;
reg_space[2135] = 8'h00;
reg_space[2136] = 8'h00;
reg_space[2137] = 8'h00;
reg_space[2138] = 8'h00;
reg_space[2139] = 8'h00;
reg_space[2140] = 8'h00;
reg_space[2141] = 8'h00;
reg_space[2142] = 8'h00;
reg_space[2143] = 8'h00;
reg_space[2144] = 8'h00;
reg_space[2145] = 8'h00;
reg_space[2146] = 8'h00;
reg_space[2147] = 8'h00;
reg_space[2148] = 8'h00;
reg_space[2149] = 8'h00;
reg_space[2150] = 8'h00;
reg_space[2151] = 8'h00;
reg_space[2152] = 8'h00;
reg_space[2153] = 8'h00;
reg_space[2154] = 8'h00;
reg_space[2155] = 8'h00;
reg_space[2156] = 8'h00;
reg_space[2157] = 8'h00;
reg_space[2158] = 8'h00;
reg_space[2159] = 8'h00;
reg_space[2160] = 8'h00;
reg_space[2161] = 8'h00;
reg_space[2162] = 8'h00;
reg_space[2163] = 8'h00;
reg_space[2164] = 8'h00;
reg_space[2165] = 8'h00;
reg_space[2166] = 8'h00;
reg_space[2167] = 8'h00;
reg_space[2168] = 8'h00;
reg_space[2169] = 8'h00;
reg_space[2170] = 8'h00;
reg_space[2171] = 8'h00;
reg_space[2172] = 8'h00;
reg_space[2173] = 8'h00;
reg_space[2174] = 8'h00;
reg_space[2175] = 8'h00;
reg_space[2176] = 8'h00;
reg_space[2177] = 8'h00;
reg_space[2178] = 8'h00;
reg_space[2179] = 8'h00;
reg_space[2180] = 8'h00;
reg_space[2181] = 8'h00;
reg_space[2182] = 8'h00;
reg_space[2183] = 8'h00;
reg_space[2184] = 8'h00;
reg_space[2185] = 8'h00;
reg_space[2186] = 8'h00;
reg_space[2187] = 8'h00;
reg_space[2188] = 8'h00;
reg_space[2189] = 8'h00;
reg_space[2190] = 8'h00;
reg_space[2191] = 8'h00;
reg_space[2192] = 8'h00;
reg_space[2193] = 8'h00;
reg_space[2194] = 8'h00;
reg_space[2195] = 8'h00;
reg_space[2196] = 8'h00;
reg_space[2197] = 8'h00;
reg_space[2198] = 8'h00;
reg_space[2199] = 8'h00;
reg_space[2200; = 8'h00;
reg_space[2201] = 8'h00;
reg_space[2202] = 8'h00;
reg_space[2203] = 8'h00;
reg_space[2204] = 8'h00;
reg_space[2205] = 8'h00;
reg_space[2206] = 8'h00;
reg_space[2207] = 8'h00;
reg_space[2208] = 8'h00;
reg_space[2209] = 8'h00;
reg_space[2210] = 8'h00;
reg_space[2211] = 8'h00;
reg_space[2212] = 8'h00;
reg_space[2213] = 8'h00;
reg_space[2214] = 8'h00;
reg_space[2215] = 8'h00;
reg_space[2216] = 8'h00;
reg_space[2217] = 8'h00;
reg_space[2218] = 8'h00;
reg_space[2219] = 8'h00;
reg_space[2220] = 8'h00;
reg_space[2221] = 8'h00;
reg_space[2222] = 8'h00;
reg_space[2223] = 8'h00;
reg_space[2224] = 8'h00;
reg_space[2225] = 8'h00;
reg_space[2226] = 8'h00;
reg_space[2227] = 8'h00;
reg_space[2228] = 8'h00;
reg_space[2229] = 8'h00;
reg_space[2230] = 8'h00;
reg_space[2231] = 8'h00;
reg_space[2232] = 8'h00;
reg_space[2233] = 8'h00;
reg_space[2234] = 8'h00;
reg_space[2235] = 8'h00;
reg_space[2236] = 8'h00;
reg_space[2237] = 8'h00;
reg_space[2238] = 8'h00;
reg_space[2239] = 8'h00;
reg_space[2240] = 8'h00;
reg_space[2241] = 8'h00;
reg_space[2242] = 8'h00;
reg_space[2243] = 8'h00;
reg_space[2244] = 8'h00;
reg_space[2245] = 8'h00;
reg_space[2246] = 8'h00;
reg_space[2247] = 8'h00;
reg_space[2248] = 8'h00;
reg_space[2249] = 8'h00;
reg_space[2250] = 8'h00;
reg_space[2251] = 8'h00;
reg_space[2252] = 8'h00;
reg_space[2253] = 8'h00;
reg_space[2254] = 8'h00;
reg_space[2255] = 8'h00;
reg_space[2256] = 8'h00;
reg_space[2257] = 8'h00;
reg_space[2258] = 8'h00;
reg_space[2259] = 8'h00;
reg_space[2260] = 8'h00;
reg_space[2261] = 8'h00;
reg_space[2262] = 8'h00;
reg_space[2263] = 8'h00;
reg_space[2264] = 8'h00;
reg_space[2265] = 8'h00;
reg_space[2266] = 8'h00;
reg_space[2267] = 8'h00;
reg_space[2268] = 8'h00;
reg_space[2269] = 8'h00;
reg_space[2270] = 8'h00;
reg_space[2271] = 8'h00;
reg_space[2272] = 8'h00;
reg_space[2273] = 8'h00;
reg_space[2274] = 8'h00;
reg_space[2275] = 8'h00;
reg_space[2276] = 8'h00;
reg_space[2277] = 8'h00;
reg_space[2278] = 8'h00;
reg_space[2279] = 8'h00;
reg_space[2280] = 8'h00;
reg_space[2281] = 8'h00;
reg_space[2282] = 8'h00;
reg_space[2283] = 8'h00;
reg_space[2284] = 8'h00;
reg_space[2285] = 8'h00;
reg_space[2286] = 8'h00;
reg_space[2287] = 8'h00;
reg_space[2288] = 8'h00;
reg_space[2289] = 8'h00;
reg_space[2290] = 8'h00;
reg_space[2291] = 8'h00;
reg_space[2292] = 8'h00;
reg_space[2293] = 8'h00;
reg_space[2294] = 8'h00;
reg_space[2295] = 8'h00;
reg_space[2296] = 8'h00;
reg_space[2297] = 8'h00;
reg_space[2298] = 8'h00;
reg_space[2299] = 8'h00;
reg_space[2300; = 8'h00;
reg_space[2301] = 8'h00;
reg_space[2302] = 8'h00;
reg_space[2303] = 8'h00;
reg_space[2304] = 8'h00;
reg_space[2305] = 8'h00;
reg_space[2306] = 8'h00;
reg_space[2307] = 8'h00;
reg_space[2308] = 8'h00;
reg_space[2309] = 8'h00;
reg_space[2310] = 8'h00;
reg_space[2311] = 8'h00;
reg_space[2312] = 8'h00;
reg_space[2313] = 8'h00;
reg_space[2314] = 8'h00;
reg_space[2315] = 8'h00;
reg_space[2316] = 8'h00;
reg_space[2317] = 8'h00;
reg_space[2318] = 8'h00;
reg_space[2319] = 8'h00;
reg_space[2320] = 8'h00;
reg_space[2321] = 8'h00;
reg_space[2322] = 8'h00;
reg_space[2323] = 8'h00;
reg_space[2324] = 8'h00;
reg_space[2325] = 8'h00;
reg_space[2326] = 8'h00;
reg_space[2327] = 8'h00;
reg_space[2328] = 8'h00;
reg_space[2329] = 8'h00;
reg_space[2330] = 8'h00;
reg_space[2331] = 8'h00;
reg_space[2332] = 8'h00;
reg_space[2333] = 8'h00;
reg_space[2334] = 8'h00;
reg_space[2335] = 8'h00;
reg_space[2336] = 8'h00;
reg_space[2337] = 8'h00;
reg_space[2338] = 8'h00;
reg_space[2339] = 8'h00;
reg_space[2340] = 8'h00;
reg_space[2341] = 8'h00;
reg_space[2342] = 8'h00;
reg_space[2343] = 8'h00;
reg_space[2344] = 8'h00;
reg_space[2345] = 8'h00;
reg_space[2346] = 8'h00;
reg_space[2347] = 8'h00;
reg_space[2348] = 8'h00;
reg_space[2349] = 8'h00;
reg_space[2350] = 8'h00;
reg_space[2351] = 8'h00;
reg_space[2352] = 8'h00;
reg_space[2353] = 8'h00;
reg_space[2354] = 8'h00;
reg_space[2355] = 8'h00;
reg_space[2356] = 8'h00;
reg_space[2357] = 8'h00;
reg_space[2358] = 8'h00;
reg_space[2359] = 8'h00;
reg_space[2360] = 8'h00;
reg_space[2361] = 8'h00;
reg_space[2362] = 8'h00;
reg_space[2363] = 8'h00;
reg_space[2364] = 8'h00;
reg_space[2365] = 8'h00;
reg_space[2366] = 8'h00;
reg_space[2367] = 8'h00;
reg_space[2368] = 8'h00;
reg_space[2369] = 8'h00;
reg_space[2370] = 8'h00;
reg_space[2371] = 8'h00;
reg_space[2372] = 8'h00;
reg_space[2373] = 8'h00;
reg_space[2374] = 8'h00;
reg_space[2375] = 8'h00;
reg_space[2376] = 8'h00;
reg_space[2377] = 8'h00;
reg_space[2378] = 8'h00;
reg_space[2379] = 8'h00;
reg_space[2380] = 8'h00;
reg_space[2381] = 8'h00;
reg_space[2382] = 8'h00;
reg_space[2383] = 8'h00;
reg_space[2384] = 8'h00;
reg_space[2385] = 8'h00;
reg_space[2386] = 8'h00;
reg_space[2387] = 8'h00;
reg_space[2388] = 8'h00;
reg_space[2389] = 8'h00;
reg_space[2390] = 8'h00;
reg_space[2391] = 8'h00;
reg_space[2392] = 8'h00;
reg_space[2393] = 8'h00;
reg_space[2394] = 8'h00;
reg_space[2395] = 8'h00;
reg_space[2396] = 8'h00;
reg_space[2397] = 8'h00;
reg_space[2398] = 8'h00;
reg_space[2399] = 8'h00;
reg_space[2400; = 8'h00;
reg_space[2401] = 8'h00;
reg_space[2402] = 8'h00;
reg_space[2403] = 8'h00;
reg_space[2404] = 8'h00;
reg_space[2405] = 8'h00;
reg_space[2406] = 8'h00;
reg_space[2407] = 8'h00;
reg_space[2408] = 8'h00;
reg_space[2409] = 8'h00;
reg_space[2410] = 8'h00;
reg_space[2411] = 8'h00;
reg_space[2412] = 8'h00;
reg_space[2413] = 8'h00;
reg_space[2414] = 8'h00;
reg_space[2415] = 8'h00;
reg_space[2416] = 8'h00;
reg_space[2417] = 8'h00;
reg_space[2418] = 8'h00;
reg_space[2419] = 8'h00;
reg_space[2420] = 8'h00;
reg_space[2421] = 8'h00;
reg_space[2422] = 8'h00;
reg_space[2423] = 8'h00;
reg_space[2424] = 8'h00;
reg_space[2425] = 8'h00;
reg_space[2426] = 8'h00;
reg_space[2427] = 8'h00;
reg_space[2428] = 8'h00;
reg_space[2429] = 8'h00;
reg_space[2430] = 8'h00;
reg_space[2431] = 8'h00;
reg_space[2432] = 8'h00;
reg_space[2433] = 8'h00;
reg_space[2434] = 8'h00;
reg_space[2435] = 8'h00;
reg_space[2436] = 8'h00;
reg_space[2437] = 8'h00;
reg_space[2438] = 8'h00;
reg_space[2439] = 8'h00;
reg_space[2440] = 8'h00;
reg_space[2441] = 8'h00;
reg_space[2442] = 8'h00;
reg_space[2443] = 8'h00;
reg_space[2444] = 8'h00;
reg_space[2445] = 8'h00;
reg_space[2446] = 8'h00;
reg_space[2447] = 8'h00;
reg_space[2448] = 8'h00;
reg_space[2449] = 8'h00;
reg_space[2450] = 8'h00;
reg_space[2451] = 8'h00;
reg_space[2452] = 8'h00;
reg_space[2453] = 8'h00;
reg_space[2454] = 8'h00;
reg_space[2455] = 8'h00;
reg_space[2456] = 8'h00;
reg_space[2457] = 8'h00;
reg_space[2458] = 8'h00;
reg_space[2459] = 8'h00;
reg_space[2460] = 8'h00;
reg_space[2461] = 8'h00;
reg_space[2462] = 8'h00;
reg_space[2463] = 8'h00;
reg_space[2464] = 8'h00;
reg_space[2465] = 8'h00;
reg_space[2466] = 8'h00;
reg_space[2467] = 8'h00;
reg_space[2468] = 8'h00;
reg_space[2469] = 8'h00;
reg_space[2470] = 8'h00;
reg_space[2471] = 8'h00;
reg_space[2472] = 8'h00;
reg_space[2473] = 8'h00;
reg_space[2474] = 8'h00;
reg_space[2475] = 8'h00;
reg_space[2476] = 8'h00;
reg_space[2477] = 8'h00;
reg_space[2478] = 8'h00;
reg_space[2479] = 8'h00;
reg_space[2480] = 8'h00;
reg_space[2481] = 8'h00;
reg_space[2482] = 8'h00;
reg_space[2483] = 8'h00;
reg_space[2484] = 8'h00;
reg_space[2485] = 8'h00;
reg_space[2486] = 8'h00;
reg_space[2487] = 8'h00;
reg_space[2488] = 8'h00;
reg_space[2489] = 8'h00;
reg_space[2490] = 8'h00;
reg_space[2491] = 8'h00;
reg_space[2492] = 8'h00;
reg_space[2493] = 8'h00;
reg_space[2494] = 8'h00;
reg_space[2495] = 8'h00;
reg_space[2496] = 8'h00;
reg_space[2497] = 8'h00;
reg_space[2498] = 8'h00;
reg_space[2499] = 8'h00;
reg_space[2500; = 8'h00;
reg_space[2501] = 8'h00;
reg_space[2502] = 8'h00;
reg_space[2503] = 8'h00;
reg_space[2504] = 8'h00;
reg_space[2505] = 8'h00;
reg_space[2506] = 8'h00;
reg_space[2507] = 8'h00;
reg_space[2508] = 8'h00;
reg_space[2509] = 8'h00;
reg_space[2510] = 8'h00;
reg_space[2511] = 8'h00;
reg_space[2512] = 8'h00;
reg_space[2513] = 8'h00;
reg_space[2514] = 8'h00;
reg_space[2515] = 8'h00;
reg_space[2516] = 8'h00;
reg_space[2517] = 8'h00;
reg_space[2518] = 8'h00;
reg_space[2519] = 8'h00;
reg_space[2520] = 8'h00;
reg_space[2521] = 8'h00;
reg_space[2522] = 8'h00;
reg_space[2523] = 8'h00;
reg_space[2524] = 8'h00;
reg_space[2525] = 8'h00;
reg_space[2526] = 8'h00;
reg_space[2527] = 8'h00;
reg_space[2528] = 8'h00;
reg_space[2529] = 8'h00;
reg_space[2530] = 8'h00;
reg_space[2531] = 8'h00;
reg_space[2532] = 8'h00;
reg_space[2533] = 8'h00;
reg_space[2534] = 8'h00;
reg_space[2535] = 8'h00;
reg_space[2536] = 8'h00;
reg_space[2537] = 8'h00;
reg_space[2538] = 8'h00;
reg_space[2539] = 8'h00;
reg_space[2540] = 8'h00;
reg_space[2541] = 8'h00;
reg_space[2542] = 8'h00;
reg_space[2543] = 8'h00;
reg_space[2544] = 8'h00;
reg_space[2545] = 8'h00;
reg_space[2546] = 8'h00;
reg_space[2547] = 8'h00;
reg_space[2548] = 8'h00;
reg_space[2549] = 8'h00;
reg_space[2550] = 8'h00;
reg_space[2551] = 8'h00;
reg_space[2552] = 8'h00;
reg_space[2553] = 8'h00;
reg_space[2554] = 8'h00;
reg_space[2555] = 8'h00;
reg_space[2556] = 8'h00;
reg_space[2557] = 8'h00;
reg_space[2558] = 8'h00;
reg_space[2559] = 8'h00;
reg_space[2560] = 8'h00;
reg_space[2561] = 8'h00;
reg_space[2562] = 8'h00;
reg_space[2563] = 8'h00;
reg_space[2564] = 8'h00;
reg_space[2565] = 8'h00;
reg_space[2566] = 8'h00;
reg_space[2567] = 8'h00;
reg_space[2568] = 8'h00;
reg_space[2569] = 8'h00;
reg_space[2570] = 8'h00;
reg_space[2571] = 8'h00;
reg_space[2572] = 8'h00;
reg_space[2573] = 8'h00;
reg_space[2574] = 8'h00;
reg_space[2575] = 8'h00;
reg_space[2576] = 8'h00;
reg_space[2577] = 8'h00;
reg_space[2578] = 8'h00;
reg_space[2579] = 8'h00;
reg_space[2580] = 8'h00;
reg_space[2581] = 8'h00;
reg_space[2582] = 8'h00;
reg_space[2583] = 8'h00;
reg_space[2584] = 8'h00;
reg_space[2585] = 8'h00;
reg_space[2586] = 8'h00;
reg_space[2587] = 8'h00;
reg_space[2588] = 8'h00;
reg_space[2589] = 8'h00;
reg_space[2590] = 8'h00;
reg_space[2591] = 8'h00;
reg_space[2592] = 8'h00;
reg_space[2593] = 8'h00;
reg_space[2594] = 8'h00;
reg_space[2595] = 8'h00;
reg_space[2596] = 8'h00;
reg_space[2597] = 8'h00;
reg_space[2598] = 8'h00;
reg_space[2599] = 8'h00;
reg_space[2600; = 8'h00;
reg_space[2601] = 8'h00;
reg_space[2602] = 8'h00;
reg_space[2603] = 8'h00;
reg_space[2604] = 8'h00;
reg_space[2605] = 8'h00;
reg_space[2606] = 8'h00;
reg_space[2607] = 8'h00;
reg_space[2608] = 8'h00;
reg_space[2609] = 8'h00;
reg_space[2610] = 8'h00;
reg_space[2611] = 8'h00;
reg_space[2612] = 8'h00;
reg_space[2613] = 8'h00;
reg_space[2614] = 8'h00;
reg_space[2615] = 8'h00;
reg_space[2616] = 8'h00;
reg_space[2617] = 8'h00;
reg_space[2618] = 8'h00;
reg_space[2619] = 8'h00;
reg_space[2620] = 8'h00;
reg_space[2621] = 8'h00;
reg_space[2622] = 8'h00;
reg_space[2623] = 8'h00;
reg_space[2624] = 8'h00;
reg_space[2625] = 8'h00;
reg_space[2626] = 8'h00;
reg_space[2627] = 8'h00;
reg_space[2628] = 8'h00;
reg_space[2629] = 8'h00;
reg_space[2630] = 8'h00;
reg_space[2631] = 8'h00;
reg_space[2632] = 8'h00;
reg_space[2633] = 8'h00;
reg_space[2634] = 8'h00;
reg_space[2635] = 8'h00;
reg_space[2636] = 8'h00;
reg_space[2637] = 8'h00;
reg_space[2638] = 8'h00;
reg_space[2639] = 8'h00;
reg_space[2640] = 8'h00;
reg_space[2641] = 8'h00;
reg_space[2642] = 8'h00;
reg_space[2643] = 8'h00;
reg_space[2644] = 8'h00;
reg_space[2645] = 8'h00;
reg_space[2646] = 8'h00;
reg_space[2647] = 8'h00;
reg_space[2648] = 8'h00;
reg_space[2649] = 8'h00;
reg_space[2650] = 8'h00;
reg_space[2651] = 8'h00;
reg_space[2652] = 8'h00;
reg_space[2653] = 8'h00;
reg_space[2654] = 8'h00;
reg_space[2655] = 8'h00;
reg_space[2656] = 8'h00;
reg_space[2657] = 8'h00;
reg_space[2658] = 8'h00;
reg_space[2659] = 8'h00;
reg_space[2660] = 8'h00;
reg_space[2661] = 8'h00;
reg_space[2662] = 8'h00;
reg_space[2663] = 8'h00;
reg_space[2664] = 8'h00;
reg_space[2665] = 8'h00;
reg_space[2666] = 8'h00;
reg_space[2667] = 8'h00;
reg_space[2668] = 8'h00;
reg_space[2669] = 8'h00;
reg_space[2670] = 8'h00;
reg_space[2671] = 8'h00;
reg_space[2672] = 8'h00;
reg_space[2673] = 8'h00;
reg_space[2674] = 8'h00;
reg_space[2675] = 8'h00;
reg_space[2676] = 8'h00;
reg_space[2677] = 8'h00;
reg_space[2678] = 8'h00;
reg_space[2679] = 8'h00;
reg_space[2680] = 8'h00;
reg_space[2681] = 8'h00;
reg_space[2682] = 8'h00;
reg_space[2683] = 8'h00;
reg_space[2684] = 8'h00;
reg_space[2685] = 8'h00;
reg_space[2686] = 8'h00;
reg_space[2687] = 8'h00;
reg_space[2688] = 8'h00;
reg_space[2689] = 8'h00;
reg_space[2690] = 8'h00;
reg_space[2691] = 8'h00;
reg_space[2692] = 8'h00;
reg_space[2693] = 8'h00;
reg_space[2694] = 8'h00;
reg_space[2695] = 8'h00;
reg_space[2696] = 8'h00;
reg_space[2697] = 8'h00;
reg_space[2698] = 8'h00;
reg_space[2699] = 8'h00;
reg_space[2700; = 8'h00;
reg_space[2701] = 8'h00;
reg_space[2702] = 8'h00;
reg_space[2703] = 8'h00;
reg_space[2704] = 8'h00;
reg_space[2705] = 8'h00;
reg_space[2706] = 8'h00;
reg_space[2707] = 8'h00;
reg_space[2708] = 8'h00;
reg_space[2709] = 8'h00;
reg_space[2710] = 8'h00;
reg_space[2711] = 8'h00;
reg_space[2712] = 8'h00;
reg_space[2713] = 8'h00;
reg_space[2714] = 8'h00;
reg_space[2715] = 8'h00;
reg_space[2716] = 8'h00;
reg_space[2717] = 8'h00;
reg_space[2718] = 8'h00;
reg_space[2719] = 8'h00;
reg_space[2720] = 8'h00;
reg_space[2721] = 8'h00;
reg_space[2722] = 8'h00;
reg_space[2723] = 8'h00;
reg_space[2724] = 8'h00;
reg_space[2725] = 8'h00;
reg_space[2726] = 8'h00;
reg_space[2727] = 8'h00;
reg_space[2728] = 8'h00;
reg_space[2729] = 8'h00;
reg_space[2730] = 8'h00;
reg_space[2731] = 8'h00;
reg_space[2732] = 8'h00;
reg_space[2733] = 8'h00;
reg_space[2734] = 8'h00;
reg_space[2735] = 8'h00;
reg_space[2736] = 8'h00;
reg_space[2737] = 8'h00;
reg_space[2738] = 8'h00;
reg_space[2739] = 8'h00;
reg_space[2740] = 8'h00;
reg_space[2741] = 8'h00;
reg_space[2742] = 8'h00;
reg_space[2743] = 8'h00;
reg_space[2744] = 8'h00;
reg_space[2745] = 8'h00;
reg_space[2746] = 8'h00;
reg_space[2747] = 8'h00;
reg_space[2748] = 8'h00;
reg_space[2749] = 8'h00;
reg_space[2750] = 8'h00;
reg_space[2751] = 8'h00;
reg_space[2752] = 8'h00;
reg_space[2753] = 8'h00;
reg_space[2754] = 8'h00;
reg_space[2755] = 8'h00;
reg_space[2756] = 8'h00;
reg_space[2757] = 8'h00;
reg_space[2758] = 8'h00;
reg_space[2759] = 8'h00;
reg_space[2760] = 8'h00;
reg_space[2761] = 8'h00;
reg_space[2762] = 8'h00;
reg_space[2763] = 8'h00;
reg_space[2764] = 8'h00;
reg_space[2765] = 8'h00;
reg_space[2766] = 8'h00;
reg_space[2767] = 8'h00;
reg_space[2768] = 8'h00;
reg_space[2769] = 8'h00;
reg_space[2770] = 8'h00;
reg_space[2771] = 8'h00;
reg_space[2772] = 8'h00;
reg_space[2773] = 8'h00;
reg_space[2774] = 8'h00;
reg_space[2775] = 8'h00;
reg_space[2776] = 8'h00;
reg_space[2777] = 8'h00;
reg_space[2778] = 8'h00;
reg_space[2779] = 8'h00;
reg_space[2780] = 8'h00;
reg_space[2781] = 8'h00;
reg_space[2782] = 8'h00;
reg_space[2783] = 8'h00;
reg_space[2784] = 8'h00;
reg_space[2785] = 8'h00;
reg_space[2786] = 8'h00;
reg_space[2787] = 8'h00;
reg_space[2788] = 8'h00;
reg_space[2789] = 8'h00;
reg_space[2790] = 8'h00;
reg_space[2791] = 8'h00;
reg_space[2792] = 8'h00;
reg_space[2793] = 8'h00;
reg_space[2794] = 8'h00;
reg_space[2795] = 8'h00;
reg_space[2796] = 8'h00;
reg_space[2797] = 8'h00;
reg_space[2798] = 8'h00;
reg_space[2799] = 8'h00;
reg_space[2800; = 8'h00;
reg_space[2801] = 8'h00;
reg_space[2802] = 8'h00;
reg_space[2803] = 8'h00;
reg_space[2804] = 8'h00;
reg_space[2805] = 8'h00;
reg_space[2806] = 8'h00;
reg_space[2807] = 8'h00;
reg_space[2808] = 8'h00;
reg_space[2809] = 8'h00;
reg_space[2810] = 8'h00;
reg_space[2811] = 8'h00;
reg_space[2812] = 8'h00;
reg_space[2813] = 8'h00;
reg_space[2814] = 8'h00;
reg_space[2815] = 8'h00;
reg_space[2816] = 8'h00;
reg_space[2817] = 8'h00;
reg_space[2818] = 8'h00;
reg_space[2819] = 8'h00;
reg_space[2820] = 8'h00;
reg_space[2821] = 8'h00;
reg_space[2822] = 8'h00;
reg_space[2823] = 8'h00;
reg_space[2824] = 8'h00;
reg_space[2825] = 8'h00;
reg_space[2826] = 8'h00;
reg_space[2827] = 8'h00;
reg_space[2828] = 8'h00;
reg_space[2829] = 8'h00;
reg_space[2830] = 8'h00;
reg_space[2831] = 8'h00;
reg_space[2832] = 8'h00;
reg_space[2833] = 8'h00;
reg_space[2834] = 8'h00;
reg_space[2835] = 8'h00;
reg_space[2836] = 8'h00;
reg_space[2837] = 8'h00;
reg_space[2838] = 8'h00;
reg_space[2839] = 8'h00;
reg_space[2840] = 8'h00;
reg_space[2841] = 8'h00;
reg_space[2842] = 8'h00;
reg_space[2843] = 8'h00;
reg_space[2844] = 8'h00;
reg_space[2845] = 8'h00;
reg_space[2846] = 8'h00;
reg_space[2847] = 8'h00;
reg_space[2848] = 8'h00;
reg_space[2849] = 8'h00;
reg_space[2850] = 8'h00;
reg_space[2851] = 8'h00;
reg_space[2852] = 8'h00;
reg_space[2853] = 8'h00;
reg_space[2854] = 8'h00;
reg_space[2855] = 8'h00;
reg_space[2856] = 8'h00;
reg_space[2857] = 8'h00;
reg_space[2858] = 8'h00;
reg_space[2859] = 8'h00;
reg_space[2860] = 8'h00;
reg_space[2861] = 8'h00;
reg_space[2862] = 8'h00;
reg_space[2863] = 8'h00;
reg_space[2864] = 8'h00;
reg_space[2865] = 8'h00;
reg_space[2866] = 8'h00;
reg_space[2867] = 8'h00;
reg_space[2868] = 8'h00;
reg_space[2869] = 8'h00;
reg_space[2870] = 8'h00;
reg_space[2871] = 8'h00;
reg_space[2872] = 8'h00;
reg_space[2873] = 8'h00;
reg_space[2874] = 8'h00;
reg_space[2875] = 8'h00;
reg_space[2876] = 8'h00;
reg_space[2877] = 8'h00;
reg_space[2878] = 8'h00;
reg_space[2879] = 8'h00;
reg_space[2880] = 8'h00;
reg_space[2881] = 8'h00;
reg_space[2882] = 8'h00;
reg_space[2883] = 8'h00;
reg_space[2884] = 8'h00;
reg_space[2885] = 8'h00;
reg_space[2886] = 8'h00;
reg_space[2887] = 8'h00;
reg_space[2888] = 8'h00;
reg_space[2889] = 8'h00;
reg_space[2890] = 8'h00;
reg_space[2891] = 8'h00;
reg_space[2892] = 8'h00;
reg_space[2893] = 8'h00;
reg_space[2894] = 8'h00;
reg_space[2895] = 8'h00;
reg_space[2896] = 8'h00;
reg_space[2897] = 8'h00;
reg_space[2898] = 8'h00;
reg_space[2899] = 8'h00;
reg_space[2900; = 8'h00;
reg_space[2901] = 8'h00;
reg_space[2902] = 8'h00;
reg_space[2903] = 8'h00;
reg_space[2904] = 8'h00;
reg_space[2905] = 8'h00;
reg_space[2906] = 8'h00;
reg_space[2907] = 8'h00;
reg_space[2908] = 8'h00;
reg_space[2909] = 8'h00;
reg_space[2910] = 8'h00;
reg_space[2911] = 8'h00;
reg_space[2912] = 8'h00;
reg_space[2913] = 8'h00;
reg_space[2914] = 8'h00;
reg_space[2915] = 8'h00;
reg_space[2916] = 8'h00;
reg_space[2917] = 8'h00;
reg_space[2918] = 8'h00;
reg_space[2919] = 8'h00;
reg_space[2920] = 8'h00;
reg_space[2921] = 8'h00;
reg_space[2922] = 8'h00;
reg_space[2923] = 8'h00;
reg_space[2924] = 8'h00;
reg_space[2925] = 8'h00;
reg_space[2926] = 8'h00;
reg_space[2927] = 8'h00;
reg_space[2928] = 8'h00;
reg_space[2929] = 8'h00;
reg_space[2930] = 8'h00;
reg_space[2931] = 8'h00;
reg_space[2932] = 8'h00;
reg_space[2933] = 8'h00;
reg_space[2934] = 8'h00;
reg_space[2935] = 8'h00;
reg_space[2936] = 8'h00;
reg_space[2937] = 8'h00;
reg_space[2938] = 8'h00;
reg_space[2939] = 8'h00;
reg_space[2940] = 8'h00;
reg_space[2941] = 8'h00;
reg_space[2942] = 8'h00;
reg_space[2943] = 8'h00;
reg_space[2944] = 8'h00;
reg_space[2945] = 8'h00;
reg_space[2946] = 8'h00;
reg_space[2947] = 8'h00;
reg_space[2948] = 8'h00;
reg_space[2949] = 8'h00;
reg_space[2950] = 8'h00;
reg_space[2951] = 8'h00;
reg_space[2952] = 8'h00;
reg_space[2953] = 8'h00;
reg_space[2954] = 8'h00;
reg_space[2955] = 8'h00;
reg_space[2956] = 8'h00;
reg_space[2957] = 8'h00;
reg_space[2958] = 8'h00;
reg_space[2959] = 8'h00;
reg_space[2960] = 8'h00;
reg_space[2961] = 8'h00;
reg_space[2962] = 8'h00;
reg_space[2963] = 8'h00;
reg_space[2964] = 8'h00;
reg_space[2965] = 8'h00;
reg_space[2966] = 8'h00;
reg_space[2967] = 8'h00;
reg_space[2968] = 8'h00;
reg_space[2969] = 8'h00;
reg_space[2970] = 8'h00;
reg_space[2971] = 8'h00;
reg_space[2972] = 8'h00;
reg_space[2973] = 8'h00;
reg_space[2974] = 8'h00;
reg_space[2975] = 8'h00;
reg_space[2976] = 8'h00;
reg_space[2977] = 8'h00;
reg_space[2978] = 8'h00;
reg_space[2979] = 8'h00;
reg_space[2980] = 8'h00;
reg_space[2981] = 8'h00;
reg_space[2982] = 8'h00;
reg_space[2983] = 8'h00;
reg_space[2984] = 8'h00;
reg_space[2985] = 8'h00;
reg_space[2986] = 8'h00;
reg_space[2987] = 8'h00;
reg_space[2988] = 8'h00;
reg_space[2989] = 8'h00;
reg_space[2990] = 8'h00;
reg_space[2991] = 8'h00;
reg_space[2992] = 8'h00;
reg_space[2993] = 8'h00;
reg_space[2994] = 8'h00;
reg_space[2995] = 8'h00;
reg_space[2996] = 8'h00;
reg_space[2997] = 8'h00;
reg_space[2998] = 8'h00;
reg_space[2999] = 8'h00;
reg_space[300;0] = 8'h00;
reg_space[300;1] = 8'h00;
reg_space[300;2] = 8'h00;
reg_space[300;3] = 8'h00;
reg_space[300;4] = 8'h00;
reg_space[300;5] = 8'h00;
reg_space[300;6] = 8'h00;
reg_space[300;7] = 8'h00;
reg_space[300;8] = 8'h00;
reg_space[300;9] = 8'h00;
reg_space[3010] = 8'h00;
reg_space[3011] = 8'h00;
reg_space[3012] = 8'h00;
reg_space[3013] = 8'h00;
reg_space[3014] = 8'h00;
reg_space[3015] = 8'h00;
reg_space[3016] = 8'h00;
reg_space[3017] = 8'h00;
reg_space[3018] = 8'h00;
reg_space[3019] = 8'h00;
reg_space[3020] = 8'h00;
reg_space[3021] = 8'h00;
reg_space[3022] = 8'h00;
reg_space[3023] = 8'h00;
reg_space[3024] = 8'h00;
reg_space[3025] = 8'h00;
reg_space[3026] = 8'h00;
reg_space[3027] = 8'h00;
reg_space[3028] = 8'h00;
reg_space[3029] = 8'h00;
reg_space[3030] = 8'h00;
reg_space[3031] = 8'h00;
reg_space[3032] = 8'h00;
reg_space[3033] = 8'h00;
reg_space[3034] = 8'h00;
reg_space[3035] = 8'h00;
reg_space[3036] = 8'h00;
reg_space[3037] = 8'h00;
reg_space[3038] = 8'h00;
reg_space[3039] = 8'h00;
reg_space[3040] = 8'h00;
reg_space[3041] = 8'h00;
reg_space[3042] = 8'h00;
reg_space[3043] = 8'h00;
reg_space[3044] = 8'h00;
reg_space[3045] = 8'h00;
reg_space[3046] = 8'h00;
reg_space[3047] = 8'h00;
reg_space[3048] = 8'h00;
reg_space[3049] = 8'h00;
reg_space[3050] = 8'h00;
reg_space[3051] = 8'h00;
reg_space[3052] = 8'h00;
reg_space[3053] = 8'h00;
reg_space[3054] = 8'h00;
reg_space[3055] = 8'h00;
reg_space[3056] = 8'h00;
reg_space[3057] = 8'h00;
reg_space[3058] = 8'h00;
reg_space[3059] = 8'h00;
reg_space[3060] = 8'h00;
reg_space[3061] = 8'h00;
reg_space[3062] = 8'h00;
reg_space[3063] = 8'h00;
reg_space[3064] = 8'h00;
reg_space[3065] = 8'h00;
reg_space[3066] = 8'h00;
reg_space[3067] = 8'h00;
reg_space[3068] = 8'h00;
reg_space[3069] = 8'h00;
reg_space[3070] = 8'h00;
reg_space[3071] = 8'h00;
reg_space[3072] = 8'h00;
reg_space[3073] = 8'h00;
reg_space[3074] = 8'h00;
reg_space[3075] = 8'h00;
reg_space[3076] = 8'h00;
reg_space[3077] = 8'h00;
reg_space[3078] = 8'h00;
reg_space[3079] = 8'h00;
reg_space[3080] = 8'h00;
reg_space[3081] = 8'h00;
reg_space[3082] = 8'h00;
reg_space[3083] = 8'h00;
reg_space[3084] = 8'h00;
reg_space[3085] = 8'h00;
reg_space[3086] = 8'h00;
reg_space[3087] = 8'h00;
reg_space[3088] = 8'h00;
reg_space[3089] = 8'h00;
reg_space[3090] = 8'h00;
reg_space[3091] = 8'h00;
reg_space[3092] = 8'h00;
reg_space[3093] = 8'h00;
reg_space[3094] = 8'h00;
reg_space[3095] = 8'h00;
reg_space[3096] = 8'h00;
reg_space[3097] = 8'h00;
reg_space[3098] = 8'h00;
reg_space[3099] = 8'h00;
reg_space[3100; = 8'h00;
reg_space[3101] = 8'h00;
reg_space[3102] = 8'h00;
reg_space[3103] = 8'h00;
reg_space[3104] = 8'h00;
reg_space[3105] = 8'h00;
reg_space[3106] = 8'h00;
reg_space[3107] = 8'h00;
reg_space[3108] = 8'h00;
reg_space[3109] = 8'h00;
reg_space[3110] = 8'h00;
reg_space[3111] = 8'h00;
reg_space[3112] = 8'h00;
reg_space[3113] = 8'h00;
reg_space[3114] = 8'h00;
reg_space[3115] = 8'h00;
reg_space[3116] = 8'h00;
reg_space[3117] = 8'h00;
reg_space[3118] = 8'h00;
reg_space[3119] = 8'h00;
reg_space[3120] = 8'h00;
reg_space[3121] = 8'h00;
reg_space[3122] = 8'h00;
reg_space[3123] = 8'h00;
reg_space[3124] = 8'h00;
reg_space[3125] = 8'h00;
reg_space[3126] = 8'h00;
reg_space[3127] = 8'h00;
reg_space[3128] = 8'h00;
reg_space[3129] = 8'h00;
reg_space[3130] = 8'h00;
reg_space[3131] = 8'h00;
reg_space[3132] = 8'h00;
reg_space[3133] = 8'h00;
reg_space[3134] = 8'h00;
reg_space[3135] = 8'h00;
reg_space[3136] = 8'h00;
reg_space[3137] = 8'h00;
reg_space[3138] = 8'h00;
reg_space[3139] = 8'h00;
reg_space[3140] = 8'h00;
reg_space[3141] = 8'h00;
reg_space[3142] = 8'h00;
reg_space[3143] = 8'h00;
reg_space[3144] = 8'h00;
reg_space[3145] = 8'h00;
reg_space[3146] = 8'h00;
reg_space[3147] = 8'h00;
reg_space[3148] = 8'h00;
reg_space[3149] = 8'h00;
reg_space[3150] = 8'h00;
reg_space[3151] = 8'h00;
reg_space[3152] = 8'h00;
reg_space[3153] = 8'h00;
reg_space[3154] = 8'h00;
reg_space[3155] = 8'h00;
reg_space[3156] = 8'h00;
reg_space[3157] = 8'h00;
reg_space[3158] = 8'h00;
reg_space[3159] = 8'h00;
reg_space[3160] = 8'h00;
reg_space[3161] = 8'h00;
reg_space[3162] = 8'h00;
reg_space[3163] = 8'h00;
reg_space[3164] = 8'h00;
reg_space[3165] = 8'h00;
reg_space[3166] = 8'h00;
reg_space[3167] = 8'h00;
reg_space[3168] = 8'h00;
reg_space[3169] = 8'h00;
reg_space[3170] = 8'h00;
reg_space[3171] = 8'h00;
reg_space[3172] = 8'h00;
reg_space[3173] = 8'h00;
reg_space[3174] = 8'h00;
reg_space[3175] = 8'h00;
reg_space[3176] = 8'h00;
reg_space[3177] = 8'h00;
reg_space[3178] = 8'h00;
reg_space[3179] = 8'h00;
reg_space[3180] = 8'h00;
reg_space[3181] = 8'h00;
reg_space[3182] = 8'h00;
reg_space[3183] = 8'h00;
reg_space[3184] = 8'h00;
reg_space[3185] = 8'h00;
reg_space[3186] = 8'h00;
reg_space[3187] = 8'h00;
reg_space[3188] = 8'h00;
reg_space[3189] = 8'h00;
reg_space[3190] = 8'h00;
reg_space[3191] = 8'h00;
reg_space[3192] = 8'h00;
reg_space[3193] = 8'h00;
reg_space[3194] = 8'h00;
reg_space[3195] = 8'h00;
reg_space[3196] = 8'h00;
reg_space[3197] = 8'h00;
reg_space[3198] = 8'h00;
reg_space[3199] = 8'h00;
reg_space[3200; = 8'h00;
reg_space[3201] = 8'h00;
reg_space[3202] = 8'h00;
reg_space[3203] = 8'h00;
reg_space[3204] = 8'h00;
reg_space[3205] = 8'h00;
reg_space[3206] = 8'h00;
reg_space[3207] = 8'h00;
reg_space[3208] = 8'h00;
reg_space[3209] = 8'h00;
reg_space[3210] = 8'h00;
reg_space[3211] = 8'h00;
reg_space[3212] = 8'h00;
reg_space[3213] = 8'h00;
reg_space[3214] = 8'h00;
reg_space[3215] = 8'h00;
reg_space[3216] = 8'h00;
reg_space[3217] = 8'h00;
reg_space[3218] = 8'h00;
reg_space[3219] = 8'h00;
reg_space[3220] = 8'h00;
reg_space[3221] = 8'h00;
reg_space[3222] = 8'h00;
reg_space[3223] = 8'h00;
reg_space[3224] = 8'h00;
reg_space[3225] = 8'h00;
reg_space[3226] = 8'h00;
reg_space[3227] = 8'h00;
reg_space[3228] = 8'h00;
reg_space[3229] = 8'h00;
reg_space[3230] = 8'h00;
reg_space[3231] = 8'h00;
reg_space[3232] = 8'h00;
reg_space[3233] = 8'h00;
reg_space[3234] = 8'h00;
reg_space[3235] = 8'h00;
reg_space[3236] = 8'h00;
reg_space[3237] = 8'h00;
reg_space[3238] = 8'h00;
reg_space[3239] = 8'h00;
reg_space[3240] = 8'h00;
reg_space[3241] = 8'h00;
reg_space[3242] = 8'h00;
reg_space[3243] = 8'h00;
reg_space[3244] = 8'h00;
reg_space[3245] = 8'h00;
reg_space[3246] = 8'h00;
reg_space[3247] = 8'h00;
reg_space[3248] = 8'h00;
reg_space[3249] = 8'h00;
reg_space[3250] = 8'h00;
reg_space[3251] = 8'h00;
reg_space[3252] = 8'h00;
reg_space[3253] = 8'h00;
reg_space[3254] = 8'h00;
reg_space[3255] = 8'h00;
reg_space[3256] = 8'h00;
reg_space[3257] = 8'h00;
reg_space[3258] = 8'h00;
reg_space[3259] = 8'h00;
reg_space[3260] = 8'h00;
reg_space[3261] = 8'h00;
reg_space[3262] = 8'h00;
reg_space[3263] = 8'h00;
reg_space[3264] = 8'h00;
reg_space[3265] = 8'h00;
reg_space[3266] = 8'h00;
reg_space[3267] = 8'h00;
reg_space[3268] = 8'h00;
reg_space[3269] = 8'h00;
reg_space[3270] = 8'h00;
reg_space[3271] = 8'h00;
reg_space[3272] = 8'h00;
reg_space[3273] = 8'h00;
reg_space[3274] = 8'h00;
reg_space[3275] = 8'h00;
reg_space[3276] = 8'h00;
reg_space[3277] = 8'h00;
reg_space[3278] = 8'h00;
reg_space[3279] = 8'h00;
reg_space[3280] = 8'h00;
reg_space[3281] = 8'h00;
reg_space[3282] = 8'h00;
reg_space[3283] = 8'h00;
reg_space[3284] = 8'h00;
reg_space[3285] = 8'h00;
reg_space[3286] = 8'h00;
reg_space[3287] = 8'h00;
reg_space[3288] = 8'h00;
reg_space[3289] = 8'h00;
reg_space[3290] = 8'h00;
reg_space[3291] = 8'h00;
reg_space[3292] = 8'h00;
reg_space[3293] = 8'h00;
reg_space[3294] = 8'h00;
reg_space[3295] = 8'h00;
reg_space[3296] = 8'h00;
reg_space[3297] = 8'h00;
reg_space[3298] = 8'h00;
reg_space[3299] = 8'h00;
reg_space[3300; = 8'h00;
reg_space[3301] = 8'h00;
reg_space[3302] = 8'h00;
reg_space[3303] = 8'h00;
reg_space[3304] = 8'h00;
reg_space[3305] = 8'h00;
reg_space[3306] = 8'h00;
reg_space[3307] = 8'h00;
reg_space[3308] = 8'h00;
reg_space[3309] = 8'h00;
reg_space[3310] = 8'h00;
reg_space[3311] = 8'h00;
reg_space[3312] = 8'h00;
reg_space[3313] = 8'h00;
reg_space[3314] = 8'h00;
reg_space[3315] = 8'h00;
reg_space[3316] = 8'h00;
reg_space[3317] = 8'h00;
reg_space[3318] = 8'h00;
reg_space[3319] = 8'h00;
reg_space[3320] = 8'h00;
reg_space[3321] = 8'h00;
reg_space[3322] = 8'h00;
reg_space[3323] = 8'h00;
reg_space[3324] = 8'h00;
reg_space[3325] = 8'h00;
reg_space[3326] = 8'h00;
reg_space[3327] = 8'h00;
reg_space[3328] = 8'h00;
reg_space[3329] = 8'h00;
reg_space[3330] = 8'h00;
reg_space[3331] = 8'h00;
reg_space[3332] = 8'h00;
reg_space[3333] = 8'h00;
reg_space[3334] = 8'h00;
reg_space[3335] = 8'h00;
reg_space[3336] = 8'h00;
reg_space[3337] = 8'h00;
reg_space[3338] = 8'h00;
reg_space[3339] = 8'h00;
reg_space[3340] = 8'h00;
reg_space[3341] = 8'h00;
reg_space[3342] = 8'h00;
reg_space[3343] = 8'h00;
reg_space[3344] = 8'h00;
reg_space[3345] = 8'h00;
reg_space[3346] = 8'h00;
reg_space[3347] = 8'h00;
reg_space[3348] = 8'h00;
reg_space[3349] = 8'h00;
reg_space[3350] = 8'h00;
reg_space[3351] = 8'h00;
reg_space[3352] = 8'h00;
reg_space[3353] = 8'h00;
reg_space[3354] = 8'h00;
reg_space[3355] = 8'h00;
reg_space[3356] = 8'h00;
reg_space[3357] = 8'h00;
reg_space[3358] = 8'h00;
reg_space[3359] = 8'h00;
reg_space[3360] = 8'h00;
reg_space[3361] = 8'h00;
reg_space[3362] = 8'h00;
reg_space[3363] = 8'h00;
reg_space[3364] = 8'h00;
reg_space[3365] = 8'h00;
reg_space[3366] = 8'h00;
reg_space[3367] = 8'h00;
reg_space[3368] = 8'h00;
reg_space[3369] = 8'h00;
reg_space[3370] = 8'h00;
reg_space[3371] = 8'h00;
reg_space[3372] = 8'h00;
reg_space[3373] = 8'h00;
reg_space[3374] = 8'h00;
reg_space[3375] = 8'h00;
reg_space[3376] = 8'h00;
reg_space[3377] = 8'h00;
reg_space[3378] = 8'h00;
reg_space[3379] = 8'h00;
reg_space[3380] = 8'h00;
reg_space[3381] = 8'h00;
reg_space[3382] = 8'h00;
reg_space[3383] = 8'h00;
reg_space[3384] = 8'h00;
reg_space[3385] = 8'h00;
reg_space[3386] = 8'h00;
reg_space[3387] = 8'h00;
reg_space[3388] = 8'h00;
reg_space[3389] = 8'h00;
reg_space[3390] = 8'h00;
reg_space[3391] = 8'h00;
reg_space[3392] = 8'h00;
reg_space[3393] = 8'h00;
reg_space[3394] = 8'h00;
reg_space[3395] = 8'h00;
reg_space[3396] = 8'h00;
reg_space[3397] = 8'h00;
reg_space[3398] = 8'h00;
reg_space[3399] = 8'h00;
reg_space[3400; = 8'h00;
reg_space[3401] = 8'h00;
reg_space[3402] = 8'h00;
reg_space[3403] = 8'h00;
reg_space[3404] = 8'h00;
reg_space[3405] = 8'h00;
reg_space[3406] = 8'h00;
reg_space[3407] = 8'h00;
reg_space[3408] = 8'h00;
reg_space[3409] = 8'h00;
reg_space[3410] = 8'h00;
reg_space[3411] = 8'h00;
reg_space[3412] = 8'h00;
reg_space[3413] = 8'h00;
reg_space[3414] = 8'h00;
reg_space[3415] = 8'h00;
reg_space[3416] = 8'h00;
reg_space[3417] = 8'h00;
reg_space[3418] = 8'h00;
reg_space[3419] = 8'h00;
reg_space[3420] = 8'h00;
reg_space[3421] = 8'h00;
reg_space[3422] = 8'h00;
reg_space[3423] = 8'h00;
reg_space[3424] = 8'h00;
reg_space[3425] = 8'h00;
reg_space[3426] = 8'h00;
reg_space[3427] = 8'h00;
reg_space[3428] = 8'h00;
reg_space[3429] = 8'h00;
reg_space[3430] = 8'h00;
reg_space[3431] = 8'h00;
reg_space[3432] = 8'h00;
reg_space[3433] = 8'h00;
reg_space[3434] = 8'h00;
reg_space[3435] = 8'h00;
reg_space[3436] = 8'h00;
reg_space[3437] = 8'h00;
reg_space[3438] = 8'h00;
reg_space[3439] = 8'h00;
reg_space[3440] = 8'h00;
reg_space[3441] = 8'h00;
reg_space[3442] = 8'h00;
reg_space[3443] = 8'h00;
reg_space[3444] = 8'h00;
reg_space[3445] = 8'h00;
reg_space[3446] = 8'h00;
reg_space[3447] = 8'h00;
reg_space[3448] = 8'h00;
reg_space[3449] = 8'h00;
reg_space[3450] = 8'h00;
reg_space[3451] = 8'h00;
reg_space[3452] = 8'h00;
reg_space[3453] = 8'h00;
reg_space[3454] = 8'h00;
reg_space[3455] = 8'h00;
reg_space[3456] = 8'h00;
reg_space[3457] = 8'h00;
reg_space[3458] = 8'h00;
reg_space[3459] = 8'h00;
reg_space[3460] = 8'h00;
reg_space[3461] = 8'h00;
reg_space[3462] = 8'h00;
reg_space[3463] = 8'h00;
reg_space[3464] = 8'h00;
reg_space[3465] = 8'h00;
reg_space[3466] = 8'h00;
reg_space[3467] = 8'h00;
reg_space[3468] = 8'h00;
reg_space[3469] = 8'h00;
reg_space[3470] = 8'h00;
reg_space[3471] = 8'h00;
reg_space[3472] = 8'h00;
reg_space[3473] = 8'h00;
reg_space[3474] = 8'h00;
reg_space[3475] = 8'h00;
reg_space[3476] = 8'h00;
reg_space[3477] = 8'h00;
reg_space[3478] = 8'h00;
reg_space[3479] = 8'h00;
reg_space[3480] = 8'h00;
reg_space[3481] = 8'h00;
reg_space[3482] = 8'h00;
reg_space[3483] = 8'h00;
reg_space[3484] = 8'h00;
reg_space[3485] = 8'h00;
reg_space[3486] = 8'h00;
reg_space[3487] = 8'h00;
reg_space[3488] = 8'h00;
reg_space[3489] = 8'h00;
reg_space[3490] = 8'h00;
reg_space[3491] = 8'h00;
reg_space[3492] = 8'h00;
reg_space[3493] = 8'h00;
reg_space[3494] = 8'h00;
reg_space[3495] = 8'h00;
reg_space[3496] = 8'h00;
reg_space[3497] = 8'h00;
reg_space[3498] = 8'h00;
reg_space[3499] = 8'h00;
reg_space[3500; = 8'h00;
reg_space[3501] = 8'h00;
reg_space[3502] = 8'h00;
reg_space[3503] = 8'h00;
reg_space[3504] = 8'h00;
reg_space[3505] = 8'h00;
reg_space[3506] = 8'h00;
reg_space[3507] = 8'h00;
reg_space[3508] = 8'h00;
reg_space[3509] = 8'h00;
reg_space[3510] = 8'h00;
reg_space[3511] = 8'h00;
reg_space[3512] = 8'h00;
reg_space[3513] = 8'h00;
reg_space[3514] = 8'h00;
reg_space[3515] = 8'h00;
reg_space[3516] = 8'h00;
reg_space[3517] = 8'h00;
reg_space[3518] = 8'h00;
reg_space[3519] = 8'h00;
reg_space[3520] = 8'h00;
reg_space[3521] = 8'h00;
reg_space[3522] = 8'h00;
reg_space[3523] = 8'h00;
reg_space[3524] = 8'h00;
reg_space[3525] = 8'h00;
reg_space[3526] = 8'h00;
reg_space[3527] = 8'h00;
reg_space[3528] = 8'h00;
reg_space[3529] = 8'h00;
reg_space[3530] = 8'h00;
reg_space[3531] = 8'h00;
reg_space[3532] = 8'h00;
reg_space[3533] = 8'h00;
reg_space[3534] = 8'h00;
reg_space[3535] = 8'h00;
reg_space[3536] = 8'h00;
reg_space[3537] = 8'h00;
reg_space[3538] = 8'h00;
reg_space[3539] = 8'h00;
reg_space[3540] = 8'h00;
reg_space[3541] = 8'h00;
reg_space[3542] = 8'h00;
reg_space[3543] = 8'h00;
reg_space[3544] = 8'h00;
reg_space[3545] = 8'h00;
reg_space[3546] = 8'h00;
reg_space[3547] = 8'h00;
reg_space[3548] = 8'h00;
reg_space[3549] = 8'h00;
reg_space[3550] = 8'h00;
reg_space[3551] = 8'h00;
reg_space[3552] = 8'h00;
reg_space[3553] = 8'h00;
reg_space[3554] = 8'h00;
reg_space[3555] = 8'h00;
reg_space[3556] = 8'h00;
reg_space[3557] = 8'h00;
reg_space[3558] = 8'h00;
reg_space[3559] = 8'h00;
reg_space[3560] = 8'h00;
reg_space[3561] = 8'h00;
reg_space[3562] = 8'h00;
reg_space[3563] = 8'h00;
reg_space[3564] = 8'h00;
reg_space[3565] = 8'h00;
reg_space[3566] = 8'h00;
reg_space[3567] = 8'h00;
reg_space[3568] = 8'h00;
reg_space[3569] = 8'h00;
reg_space[3570] = 8'h00;
reg_space[3571] = 8'h00;
reg_space[3572] = 8'h00;
reg_space[3573] = 8'h00;
reg_space[3574] = 8'h00;
reg_space[3575] = 8'h00;
reg_space[3576] = 8'h00;
reg_space[3577] = 8'h00;
reg_space[3578] = 8'h00;
reg_space[3579] = 8'h00;
reg_space[3580] = 8'h00;
reg_space[3581] = 8'h00;
reg_space[3582] = 8'h00;
reg_space[3583] = 8'h00;
reg_space[3584] = 8'h00;
reg_space[3585] = 8'h00;
reg_space[3586] = 8'h00;
reg_space[3587] = 8'h00;
reg_space[3588] = 8'h00;
reg_space[3589] = 8'h00;
reg_space[3590] = 8'h00;
reg_space[3591] = 8'h00;
reg_space[3592] = 8'h00;
reg_space[3593] = 8'h00;
reg_space[3594] = 8'h00;
reg_space[3595] = 8'h00;
reg_space[3596] = 8'h00;
reg_space[3597] = 8'h00;
reg_space[3598] = 8'h00;
reg_space[3599] = 8'h00;
reg_space[3600; = 8'h00;
reg_space[3601] = 8'h00;
reg_space[3602] = 8'h00;
reg_space[3603] = 8'h00;
reg_space[3604] = 8'h00;
reg_space[3605] = 8'h00;
reg_space[3606] = 8'h00;
reg_space[3607] = 8'h00;
reg_space[3608] = 8'h00;
reg_space[3609] = 8'h00;
reg_space[3610] = 8'h00;
reg_space[3611] = 8'h00;
reg_space[3612] = 8'h00;
reg_space[3613] = 8'h00;
reg_space[3614] = 8'h00;
reg_space[3615] = 8'h00;
reg_space[3616] = 8'h00;
reg_space[3617] = 8'h00;
reg_space[3618] = 8'h00;
reg_space[3619] = 8'h00;
reg_space[3620] = 8'h00;
reg_space[3621] = 8'h00;
reg_space[3622] = 8'h00;
reg_space[3623] = 8'h00;
reg_space[3624] = 8'h00;
reg_space[3625] = 8'h00;
reg_space[3626] = 8'h00;
reg_space[3627] = 8'h00;
reg_space[3628] = 8'h00;
reg_space[3629] = 8'h00;
reg_space[3630] = 8'h00;
reg_space[3631] = 8'h00;
reg_space[3632] = 8'h00;
reg_space[3633] = 8'h00;
reg_space[3634] = 8'h00;
reg_space[3635] = 8'h00;
reg_space[3636] = 8'h00;
reg_space[3637] = 8'h00;
reg_space[3638] = 8'h00;
reg_space[3639] = 8'h00;
reg_space[3640] = 8'h00;
reg_space[3641] = 8'h00;
reg_space[3642] = 8'h00;
reg_space[3643] = 8'h00;
reg_space[3644] = 8'h00;
reg_space[3645] = 8'h00;
reg_space[3646] = 8'h00;
reg_space[3647] = 8'h00;
reg_space[3648] = 8'h00;
reg_space[3649] = 8'h00;
reg_space[3650] = 8'h00;
reg_space[3651] = 8'h00;
reg_space[3652] = 8'h00;
reg_space[3653] = 8'h00;
reg_space[3654] = 8'h00;
reg_space[3655] = 8'h00;
reg_space[3656] = 8'h00;
reg_space[3657] = 8'h00;
reg_space[3658] = 8'h00;
reg_space[3659] = 8'h00;
reg_space[3660] = 8'h00;
reg_space[3661] = 8'h00;
reg_space[3662] = 8'h00;
reg_space[3663] = 8'h00;
reg_space[3664] = 8'h00;
reg_space[3665] = 8'h00;
reg_space[3666] = 8'h00;
reg_space[3667] = 8'h00;
reg_space[3668] = 8'h00;
reg_space[3669] = 8'h00;
reg_space[3670] = 8'h00;
reg_space[3671] = 8'h00;
reg_space[3672] = 8'h00;
reg_space[3673] = 8'h00;
reg_space[3674] = 8'h00;
reg_space[3675] = 8'h00;
reg_space[3676] = 8'h00;
reg_space[3677] = 8'h00;
reg_space[3678] = 8'h00;
reg_space[3679] = 8'h00;
reg_space[3680] = 8'h00;
reg_space[3681] = 8'h00;
reg_space[3682] = 8'h00;
reg_space[3683] = 8'h00;
reg_space[3684] = 8'h00;
reg_space[3685] = 8'h00;
reg_space[3686] = 8'h00;
reg_space[3687] = 8'h00;
reg_space[3688] = 8'h00;
reg_space[3689] = 8'h00;
reg_space[3690] = 8'h00;
reg_space[3691] = 8'h00;
reg_space[3692] = 8'h00;
reg_space[3693] = 8'h00;
reg_space[3694] = 8'h00;
reg_space[3695] = 8'h00;
reg_space[3696] = 8'h00;
reg_space[3697] = 8'h00;
reg_space[3698] = 8'h00;
reg_space[3699] = 8'h00;
reg_space[3700; = 8'h00;
reg_space[3701] = 8'h00;
reg_space[3702] = 8'h00;
reg_space[3703] = 8'h00;
reg_space[3704] = 8'h00;
reg_space[3705] = 8'h00;
reg_space[3706] = 8'h00;
reg_space[3707] = 8'h00;
reg_space[3708] = 8'h00;
reg_space[3709] = 8'h00;
reg_space[3710] = 8'h00;
reg_space[3711] = 8'h00;
reg_space[3712] = 8'h00;
reg_space[3713] = 8'h00;
reg_space[3714] = 8'h00;
reg_space[3715] = 8'h00;
reg_space[3716] = 8'h00;
reg_space[3717] = 8'h00;
reg_space[3718] = 8'h00;
reg_space[3719] = 8'h00;
reg_space[3720] = 8'h00;
reg_space[3721] = 8'h00;
reg_space[3722] = 8'h00;
reg_space[3723] = 8'h00;
reg_space[3724] = 8'h00;
reg_space[3725] = 8'h00;
reg_space[3726] = 8'h00;
reg_space[3727] = 8'h00;
reg_space[3728] = 8'h00;
reg_space[3729] = 8'h00;
reg_space[3730] = 8'h00;
reg_space[3731] = 8'h00;
reg_space[3732] = 8'h00;
reg_space[3733] = 8'h00;
reg_space[3734] = 8'h00;
reg_space[3735] = 8'h00;
reg_space[3736] = 8'h00;
reg_space[3737] = 8'h00;
reg_space[3738] = 8'h00;
reg_space[3739] = 8'h00;
reg_space[3740] = 8'h00;
reg_space[3741] = 8'h00;
reg_space[3742] = 8'h00;
reg_space[3743] = 8'h00;
reg_space[3744] = 8'h00;
reg_space[3745] = 8'h00;
reg_space[3746] = 8'h00;
reg_space[3747] = 8'h00;
reg_space[3748] = 8'h00;
reg_space[3749] = 8'h00;
reg_space[3750] = 8'h00;
reg_space[3751] = 8'h00;
reg_space[3752] = 8'h00;
reg_space[3753] = 8'h00;
reg_space[3754] = 8'h00;
reg_space[3755] = 8'h00;
reg_space[3756] = 8'h00;
reg_space[3757] = 8'h00;
reg_space[3758] = 8'h00;
reg_space[3759] = 8'h00;
reg_space[3760] = 8'h00;
reg_space[3761] = 8'h00;
reg_space[3762] = 8'h00;
reg_space[3763] = 8'h00;
reg_space[3764] = 8'h00;
reg_space[3765] = 8'h00;
reg_space[3766] = 8'h00;
reg_space[3767] = 8'h00;
reg_space[3768] = 8'h00;
reg_space[3769] = 8'h00;
reg_space[3770] = 8'h00;
reg_space[3771] = 8'h00;
reg_space[3772] = 8'h00;
reg_space[3773] = 8'h00;
reg_space[3774] = 8'h00;
reg_space[3775] = 8'h00;
reg_space[3776] = 8'h00;
reg_space[3777] = 8'h00;
reg_space[3778] = 8'h00;
reg_space[3779] = 8'h00;
reg_space[3780] = 8'h00;
reg_space[3781] = 8'h00;
reg_space[3782] = 8'h00;
reg_space[3783] = 8'h00;
reg_space[3784] = 8'h00;
reg_space[3785] = 8'h00;
reg_space[3786] = 8'h00;
reg_space[3787] = 8'h00;
reg_space[3788] = 8'h00;
reg_space[3789] = 8'h00;
reg_space[3790] = 8'h00;
reg_space[3791] = 8'h00;
reg_space[3792] = 8'h00;
reg_space[3793] = 8'h00;
reg_space[3794] = 8'h00;
reg_space[3795] = 8'h00;
reg_space[3796] = 8'h00;
reg_space[3797] = 8'h00;
reg_space[3798] = 8'h00;
reg_space[3799] = 8'h00;
reg_space[3800; = 8'h00;
reg_space[3801] = 8'h00;
reg_space[3802] = 8'h00;
reg_space[3803] = 8'h00;
reg_space[3804] = 8'h00;
reg_space[3805] = 8'h00;
reg_space[3806] = 8'h00;
reg_space[3807] = 8'h00;
reg_space[3808] = 8'h00;
reg_space[3809] = 8'h00;
reg_space[3810] = 8'h00;
reg_space[3811] = 8'h00;
reg_space[3812] = 8'h00;
reg_space[3813] = 8'h00;
reg_space[3814] = 8'h00;
reg_space[3815] = 8'h00;
reg_space[3816] = 8'h00;
reg_space[3817] = 8'h00;
reg_space[3818] = 8'h00;
reg_space[3819] = 8'h00;
reg_space[3820] = 8'h00;
reg_space[3821] = 8'h00;
reg_space[3822] = 8'h00;
reg_space[3823] = 8'h00;
reg_space[3824] = 8'h00;
reg_space[3825] = 8'h00;
reg_space[3826] = 8'h00;
reg_space[3827] = 8'h00;
reg_space[3828] = 8'h00;
reg_space[3829] = 8'h00;
reg_space[3830] = 8'h00;
reg_space[3831] = 8'h00;
reg_space[3832] = 8'h00;
reg_space[3833] = 8'h00;
reg_space[3834] = 8'h00;
reg_space[3835] = 8'h00;
reg_space[3836] = 8'h00;
reg_space[3837] = 8'h00;
reg_space[3838] = 8'h00;
reg_space[3839] = 8'h00;
reg_space[3840] = 8'h00;
reg_space[3841] = 8'h00;
reg_space[3842] = 8'h00;
reg_space[3843] = 8'h00;
reg_space[3844] = 8'h00;
reg_space[3845] = 8'h00;
reg_space[3846] = 8'h00;
reg_space[3847] = 8'h00;
reg_space[3848] = 8'h00;
reg_space[3849] = 8'h00;
reg_space[3850] = 8'h00;
reg_space[3851] = 8'h00;
reg_space[3852] = 8'h00;
reg_space[3853] = 8'h00;
reg_space[3854] = 8'h00;
reg_space[3855] = 8'h00;
reg_space[3856] = 8'h00;
reg_space[3857] = 8'h00;
reg_space[3858] = 8'h00;
reg_space[3859] = 8'h00;
reg_space[3860] = 8'h00;
reg_space[3861] = 8'h00;
reg_space[3862] = 8'h00;
reg_space[3863] = 8'h00;
reg_space[3864] = 8'h00;
reg_space[3865] = 8'h00;
reg_space[3866] = 8'h00;
reg_space[3867] = 8'h00;
reg_space[3868] = 8'h00;
reg_space[3869] = 8'h00;
reg_space[3870] = 8'h00;
reg_space[3871] = 8'h00;
reg_space[3872] = 8'h00;
reg_space[3873] = 8'h00;
reg_space[3874] = 8'h00;
reg_space[3875] = 8'h00;
reg_space[3876] = 8'h00;
reg_space[3877] = 8'h00;
reg_space[3878] = 8'h00;
reg_space[3879] = 8'h00;
reg_space[3880] = 8'h00;
reg_space[3881] = 8'h00;
reg_space[3882] = 8'h00;
reg_space[3883] = 8'h00;
reg_space[3884] = 8'h00;
reg_space[3885] = 8'h00;
reg_space[3886] = 8'h00;
reg_space[3887] = 8'h00;
reg_space[3888] = 8'h00;
reg_space[3889] = 8'h00;
reg_space[3890] = 8'h00;
reg_space[3891] = 8'h00;
reg_space[3892] = 8'h00;
reg_space[3893] = 8'h00;
reg_space[3894] = 8'h00;
reg_space[3895] = 8'h00;
reg_space[3896] = 8'h00;
reg_space[3897] = 8'h00;
reg_space[3898] = 8'h00;
reg_space[3899] = 8'h00;
reg_space[3900; = 8'h00;
reg_space[3901] = 8'h00;
reg_space[3902] = 8'h00;
reg_space[3903] = 8'h00;
reg_space[3904] = 8'h00;
reg_space[3905] = 8'h00;
reg_space[3906] = 8'h00;
reg_space[3907] = 8'h00;
reg_space[3908] = 8'h00;
reg_space[3909] = 8'h00;
reg_space[3910] = 8'h00;
reg_space[3911] = 8'h00;
reg_space[3912] = 8'h00;
reg_space[3913] = 8'h00;
reg_space[3914] = 8'h00;
reg_space[3915] = 8'h00;
reg_space[3916] = 8'h00;
reg_space[3917] = 8'h00;
reg_space[3918] = 8'h00;
reg_space[3919] = 8'h00;
reg_space[3920] = 8'h00;
reg_space[3921] = 8'h00;
reg_space[3922] = 8'h00;
reg_space[3923] = 8'h00;
reg_space[3924] = 8'h00;
reg_space[3925] = 8'h00;
reg_space[3926] = 8'h00;
reg_space[3927] = 8'h00;
reg_space[3928] = 8'h00;
reg_space[3929] = 8'h00;
reg_space[3930] = 8'h00;
reg_space[3931] = 8'h00;
reg_space[3932] = 8'h00;
reg_space[3933] = 8'h00;
reg_space[3934] = 8'h00;
reg_space[3935] = 8'h00;
reg_space[3936] = 8'h00;
reg_space[3937] = 8'h00;
reg_space[3938] = 8'h00;
reg_space[3939] = 8'h00;
reg_space[3940] = 8'h00;
reg_space[3941] = 8'h00;
reg_space[3942] = 8'h00;
reg_space[3943] = 8'h00;
reg_space[3944] = 8'h00;
reg_space[3945] = 8'h00;
reg_space[3946] = 8'h00;
reg_space[3947] = 8'h00;
reg_space[3948] = 8'h00;
reg_space[3949] = 8'h00;
reg_space[3950] = 8'h00;
reg_space[3951] = 8'h00;
reg_space[3952] = 8'h00;
reg_space[3953] = 8'h00;
reg_space[3954] = 8'h00;
reg_space[3955] = 8'h00;
reg_space[3956] = 8'h00;
reg_space[3957] = 8'h00;
reg_space[3958] = 8'h00;
reg_space[3959] = 8'h00;
reg_space[3960] = 8'h00;
reg_space[3961] = 8'h00;
reg_space[3962] = 8'h00;
reg_space[3963] = 8'h00;
reg_space[3964] = 8'h00;
reg_space[3965] = 8'h00;
reg_space[3966] = 8'h00;
reg_space[3967] = 8'h00;
reg_space[3968] = 8'h00;
reg_space[3969] = 8'h00;
reg_space[3970] = 8'h00;
reg_space[3971] = 8'h00;
reg_space[3972] = 8'h00;
reg_space[3973] = 8'h00;
reg_space[3974] = 8'h00;
reg_space[3975] = 8'h00;
reg_space[3976] = 8'h00;
reg_space[3977] = 8'h00;
reg_space[3978] = 8'h00;
reg_space[3979] = 8'h00;
reg_space[3980] = 8'h00;
reg_space[3981] = 8'h00;
reg_space[3982] = 8'h00;
reg_space[3983] = 8'h00;
reg_space[3984] = 8'h00;
reg_space[3985] = 8'h00;
reg_space[3986] = 8'h00;
reg_space[3987] = 8'h00;
reg_space[3988] = 8'h00;
reg_space[3989] = 8'h00;
reg_space[3990] = 8'h00;
reg_space[3991] = 8'h00;
reg_space[3992] = 8'h00;
reg_space[3993] = 8'h00;
reg_space[3994] = 8'h00;
reg_space[3995] = 8'h00;
reg_space[3996] = 8'h00;
reg_space[3997] = 8'h00;
reg_space[3998] = 8'h00;
reg_space[3999] = 8'h00;
reg_space[400;0] = 8'h00;
reg_space[400;1] = 8'h00;
reg_space[400;2] = 8'h00;
reg_space[400;3] = 8'h00;
reg_space[400;4] = 8'h00;
reg_space[400;5] = 8'h00;
reg_space[400;6] = 8'h00;
reg_space[400;7] = 8'h00;
reg_space[400;8] = 8'h00;
reg_space[400;9] = 8'h00;
reg_space[4010] = 8'h00;
reg_space[4011] = 8'h00;
reg_space[4012] = 8'h00;
reg_space[4013] = 8'h00;
reg_space[4014] = 8'h00;
reg_space[4015] = 8'h00;
reg_space[4016] = 8'h00;
reg_space[4017] = 8'h00;
reg_space[4018] = 8'h00;
reg_space[4019] = 8'h00;
reg_space[4020] = 8'h00;
reg_space[4021] = 8'h00;
reg_space[4022] = 8'h00;
reg_space[4023] = 8'h00;
reg_space[4024] = 8'h00;
reg_space[4025] = 8'h00;
reg_space[4026] = 8'h00;
reg_space[4027] = 8'h00;
reg_space[4028] = 8'h00;
reg_space[4029] = 8'h00;
reg_space[4030] = 8'h00;
reg_space[4031] = 8'h00;
reg_space[4032] = 8'h00;
reg_space[4033] = 8'h00;
reg_space[4034] = 8'h00;
reg_space[4035] = 8'h00;
reg_space[4036] = 8'h00;
reg_space[4037] = 8'h00;
reg_space[4038] = 8'h00;
reg_space[4039] = 8'h00;
reg_space[4040] = 8'h00;
reg_space[4041] = 8'h00;
reg_space[4042] = 8'h00;
reg_space[4043] = 8'h00;
reg_space[4044] = 8'h00;
reg_space[4045] = 8'h00;
reg_space[4046] = 8'h00;
reg_space[4047] = 8'h00;
reg_space[4048] = 8'h00;
reg_space[4049] = 8'h00;
reg_space[4050] = 8'h00;
reg_space[4051] = 8'h00;
reg_space[4052] = 8'h00;
reg_space[4053] = 8'h00;
reg_space[4054] = 8'h00;
reg_space[4055] = 8'h00;
reg_space[4056] = 8'h00;
reg_space[4057] = 8'h00;
reg_space[4058] = 8'h00;
reg_space[4059] = 8'h00;
reg_space[4060] = 8'h00;
reg_space[4061] = 8'h00;
reg_space[4062] = 8'h00;
reg_space[4063] = 8'h00;
reg_space[4064] = 8'h00;
reg_space[4065] = 8'h00;
reg_space[4066] = 8'h00;
reg_space[4067] = 8'h00;
reg_space[4068] = 8'h00;
reg_space[4069] = 8'h00;
reg_space[4070] = 8'h00;
reg_space[4071] = 8'h00;
reg_space[4072] = 8'h00;
reg_space[4073] = 8'h00;
reg_space[4074] = 8'h00;
reg_space[4075] = 8'h00;
reg_space[4076] = 8'h00;
reg_space[4077] = 8'h00;
reg_space[4078] = 8'h00;
reg_space[4079] = 8'h00;
reg_space[4080] = 8'h00;
reg_space[4081] = 8'h00;
reg_space[4082] = 8'h00;
reg_space[4083] = 8'h00;
reg_space[4084] = 8'h00;
reg_space[4085] = 8'h00;
reg_space[4086] = 8'h00;
reg_space[4087] = 8'h00;
reg_space[4088] = 8'h00;
reg_space[4089] = 8'h00;
reg_space[4090] = 8'h00;
reg_space[4091] = 8'h00;
reg_space[4092] = 8'h00;
reg_space[4093] = 8'h00;
reg_space[4094] = 8'h00;
reg_space[4095] = 8'h00;
reg_space[4096] = 8'h00;
reg_space[4097] = 8'h00;
reg_space[4098] = 8'h00;
reg_space[4099] = 8'h00;
reg_space[4100; = 8'h00;
reg_space[4101] = 8'h00;
reg_space[4102] = 8'h00;
reg_space[4103] = 8'h00;
reg_space[4104] = 8'h00;
reg_space[4105] = 8'h00;
reg_space[4106] = 8'h00;
reg_space[4107] = 8'h00;
reg_space[4108] = 8'h00;
reg_space[4109] = 8'h00;
reg_space[4110] = 8'h00;
reg_space[4111] = 8'h00;
reg_space[4112] = 8'h00;
reg_space[4113] = 8'h00;
reg_space[4114] = 8'h00;
reg_space[4115] = 8'h00;
reg_space[4116] = 8'h00;
reg_space[4117] = 8'h00;
reg_space[4118] = 8'h00;
reg_space[4119] = 8'h00;
reg_space[4120] = 8'h00;
reg_space[4121] = 8'h00;
reg_space[4122] = 8'h00;
reg_space[4123] = 8'h00;
reg_space[4124] = 8'h00;
reg_space[4125] = 8'h00;
reg_space[4126] = 8'h00;
reg_space[4127] = 8'h00;
reg_space[4128] = 8'h00;
reg_space[4129] = 8'h00;
reg_space[4130] = 8'h00;
reg_space[4131] = 8'h00;
reg_space[4132] = 8'h00;
reg_space[4133] = 8'h00;
reg_space[4134] = 8'h00;
reg_space[4135] = 8'h00;
reg_space[4136] = 8'h00;
reg_space[4137] = 8'h00;
reg_space[4138] = 8'h00;
reg_space[4139] = 8'h00;
reg_space[4140] = 8'h00;
reg_space[4141] = 8'h00;
reg_space[4142] = 8'h00;
reg_space[4143] = 8'h00;
reg_space[4144] = 8'h00;
reg_space[4145] = 8'h00;
reg_space[4146] = 8'h00;
reg_space[4147] = 8'h00;
reg_space[4148] = 8'h00;
reg_space[4149] = 8'h00;
reg_space[4150] = 8'h00;
reg_space[4151] = 8'h00;
reg_space[4152] = 8'h00;
reg_space[4153] = 8'h00;
reg_space[4154] = 8'h00;
reg_space[4155] = 8'h00;
reg_space[4156] = 8'h00;
reg_space[4157] = 8'h00;
reg_space[4158] = 8'h00;
reg_space[4159] = 8'h00;
reg_space[4160] = 8'h00;
reg_space[4161] = 8'h00;
reg_space[4162] = 8'h00;
reg_space[4163] = 8'h00;
reg_space[4164] = 8'h00;
reg_space[4165] = 8'h00;
reg_space[4166] = 8'h00;
reg_space[4167] = 8'h00;
reg_space[4168] = 8'h00;
reg_space[4169] = 8'h00;
reg_space[4170] = 8'h00;
reg_space[4171] = 8'h00;
reg_space[4172] = 8'h00;
reg_space[4173] = 8'h00;
reg_space[4174] = 8'h00;
reg_space[4175] = 8'h00;
reg_space[4176] = 8'h00;
reg_space[4177] = 8'h00;
reg_space[4178] = 8'h00;
reg_space[4179] = 8'h00;
reg_space[4180] = 8'h00;
reg_space[4181] = 8'h00;
reg_space[4182] = 8'h00;
reg_space[4183] = 8'h00;
reg_space[4184] = 8'h00;
reg_space[4185] = 8'h00;
reg_space[4186] = 8'h00;
reg_space[4187] = 8'h00;
reg_space[4188] = 8'h00;
reg_space[4189] = 8'h00;
reg_space[4190] = 8'h00;
reg_space[4191] = 8'h00;
reg_space[4192] = 8'h00;
reg_space[4193] = 8'h00;
reg_space[4194] = 8'h00;
reg_space[4195] = 8'h00;
reg_space[4196] = 8'h00;
reg_space[4197] = 8'h00;
reg_space[4198] = 8'h00;
reg_space[4199] = 8'h00;
reg_space[4200; = 8'h00;
reg_space[4201] = 8'h00;
reg_space[4202] = 8'h00;
reg_space[4203] = 8'h00;
reg_space[4204] = 8'h00;
reg_space[4205] = 8'h00;
reg_space[4206] = 8'h00;
reg_space[4207] = 8'h00;
reg_space[4208] = 8'h00;
reg_space[4209] = 8'h00;
reg_space[4210] = 8'h00;
reg_space[4211] = 8'h00;
reg_space[4212] = 8'h00;
reg_space[4213] = 8'h00;
reg_space[4214] = 8'h00;
reg_space[4215] = 8'h00;
reg_space[4216] = 8'h00;
reg_space[4217] = 8'h00;
reg_space[4218] = 8'h00;
reg_space[4219] = 8'h00;
reg_space[4220] = 8'h00;
reg_space[4221] = 8'h00;
reg_space[4222] = 8'h00;
reg_space[4223] = 8'h00;
reg_space[4224] = 8'h00;
reg_space[4225] = 8'h00;
reg_space[4226] = 8'h00;
reg_space[4227] = 8'h00;
reg_space[4228] = 8'h00;
reg_space[4229] = 8'h00;
reg_space[4230] = 8'h00;
reg_space[4231] = 8'h00;
reg_space[4232] = 8'h00;
reg_space[4233] = 8'h00;
reg_space[4234] = 8'h00;
reg_space[4235] = 8'h00;
reg_space[4236] = 8'h00;
reg_space[4237] = 8'h00;
reg_space[4238] = 8'h00;
reg_space[4239] = 8'h00;
reg_space[4240] = 8'h00;
reg_space[4241] = 8'h00;
reg_space[4242] = 8'h00;
reg_space[4243] = 8'h00;
reg_space[4244] = 8'h00;
reg_space[4245] = 8'h00;
reg_space[4246] = 8'h00;
reg_space[4247] = 8'h00;
reg_space[4248] = 8'h00;
reg_space[4249] = 8'h00;
reg_space[4250] = 8'h00;
reg_space[4251] = 8'h00;
reg_space[4252] = 8'h00;
reg_space[4253] = 8'h00;
reg_space[4254] = 8'h00;
reg_space[4255] = 8'h00;
reg_space[4256] = 8'h00;
reg_space[4257] = 8'h00;
reg_space[4258] = 8'h00;
reg_space[4259] = 8'h00;
reg_space[4260] = 8'h00;
reg_space[4261] = 8'h00;
reg_space[4262] = 8'h00;
reg_space[4263] = 8'h00;
reg_space[4264] = 8'h00;
reg_space[4265] = 8'h00;
reg_space[4266] = 8'h00;
reg_space[4267] = 8'h00;
reg_space[4268] = 8'h00;
reg_space[4269] = 8'h00;
reg_space[4270] = 8'h00;
reg_space[4271] = 8'h00;
reg_space[4272] = 8'h00;
reg_space[4273] = 8'h00;
reg_space[4274] = 8'h00;
reg_space[4275] = 8'h00;
reg_space[4276] = 8'h00;
reg_space[4277] = 8'h00;
reg_space[4278] = 8'h00;
reg_space[4279] = 8'h00;
reg_space[4280] = 8'h00;
reg_space[4281] = 8'h00;
reg_space[4282] = 8'h00;
reg_space[4283] = 8'h00;
reg_space[4284] = 8'h00;
reg_space[4285] = 8'h00;
reg_space[4286] = 8'h00;
reg_space[4287] = 8'h00;
reg_space[4288] = 8'h00;
reg_space[4289] = 8'h00;
reg_space[4290] = 8'h00;
reg_space[4291] = 8'h00;
reg_space[4292] = 8'h00;
reg_space[4293] = 8'h00;
reg_space[4294] = 8'h00;
reg_space[4295] = 8'h00;
reg_space[4296] = 8'h00;
reg_space[4297] = 8'h00;
reg_space[4298] = 8'h00;
reg_space[4299] = 8'h00;
reg_space[4300; = 8'h00;
reg_space[4301] = 8'h00;
reg_space[4302] = 8'h00;
reg_space[4303] = 8'h00;
reg_space[4304] = 8'h00;
reg_space[4305] = 8'h00;
reg_space[4306] = 8'h00;
reg_space[4307] = 8'h00;
reg_space[4308] = 8'h00;
reg_space[4309] = 8'h00;
reg_space[4310] = 8'h00;
reg_space[4311] = 8'h00;
reg_space[4312] = 8'h00;
reg_space[4313] = 8'h00;
reg_space[4314] = 8'h00;
reg_space[4315] = 8'h00;
reg_space[4316] = 8'h00;
reg_space[4317] = 8'h00;
reg_space[4318] = 8'h00;
reg_space[4319] = 8'h00;
reg_space[4320] = 8'h00;
reg_space[4321] = 8'h00;
reg_space[4322] = 8'h00;
reg_space[4323] = 8'h00;
reg_space[4324] = 8'h00;
reg_space[4325] = 8'h00;
reg_space[4326] = 8'h00;
reg_space[4327] = 8'h00;
reg_space[4328] = 8'h00;
reg_space[4329] = 8'h00;
reg_space[4330] = 8'h00;
reg_space[4331] = 8'h00;
reg_space[4332] = 8'h00;
reg_space[4333] = 8'h00;
reg_space[4334] = 8'h00;
reg_space[4335] = 8'h00;
reg_space[4336] = 8'h00;
reg_space[4337] = 8'h00;
reg_space[4338] = 8'h00;
reg_space[4339] = 8'h00;
reg_space[4340] = 8'h00;
reg_space[4341] = 8'h00;
reg_space[4342] = 8'h00;
reg_space[4343] = 8'h00;
reg_space[4344] = 8'h00;
reg_space[4345] = 8'h00;
reg_space[4346] = 8'h00;
reg_space[4347] = 8'h00;
reg_space[4348] = 8'h00;
reg_space[4349] = 8'h00;
reg_space[4350] = 8'h00;
reg_space[4351] = 8'h00;
reg_space[4352] = 8'h00;
reg_space[4353] = 8'h00;
reg_space[4354] = 8'h00;
reg_space[4355] = 8'h00;
reg_space[4356] = 8'h00;
reg_space[4357] = 8'h00;
reg_space[4358] = 8'h00;
reg_space[4359] = 8'h00;
reg_space[4360] = 8'h00;
reg_space[4361] = 8'h00;
reg_space[4362] = 8'h00;
reg_space[4363] = 8'h00;
reg_space[4364] = 8'h00;
reg_space[4365] = 8'h00;
reg_space[4366] = 8'h00;
reg_space[4367] = 8'h00;
reg_space[4368] = 8'h00;
reg_space[4369] = 8'h00;
reg_space[4370] = 8'h00;
reg_space[4371] = 8'h00;
reg_space[4372] = 8'h00;
reg_space[4373] = 8'h00;
reg_space[4374] = 8'h00;
reg_space[4375] = 8'h00;
reg_space[4376] = 8'h00;
reg_space[4377] = 8'h00;
reg_space[4378] = 8'h00;
reg_space[4379] = 8'h00;
reg_space[4380] = 8'h00;
reg_space[4381] = 8'h00;
reg_space[4382] = 8'h00;
reg_space[4383] = 8'h00;
reg_space[4384] = 8'h00;
reg_space[4385] = 8'h00;
reg_space[4386] = 8'h00;
reg_space[4387] = 8'h00;
reg_space[4388] = 8'h00;
reg_space[4389] = 8'h00;
reg_space[4390] = 8'h00;
reg_space[4391] = 8'h00;
reg_space[4392] = 8'h00;
reg_space[4393] = 8'h00;
reg_space[4394] = 8'h00;
reg_space[4395] = 8'h00;
reg_space[4396] = 8'h00;
reg_space[4397] = 8'h00;
reg_space[4398] = 8'h00;
reg_space[4399] = 8'h00;
reg_space[4400; = 8'h00;
reg_space[4401] = 8'h00;
reg_space[4402] = 8'h00;
reg_space[4403] = 8'h00;
reg_space[4404] = 8'h00;
reg_space[4405] = 8'h00;
reg_space[4406] = 8'h00;
reg_space[4407] = 8'h00;
reg_space[4408] = 8'h00;
reg_space[4409] = 8'h00;
reg_space[4410] = 8'h00;
reg_space[4411] = 8'h00;
reg_space[4412] = 8'h00;
reg_space[4413] = 8'h00;
reg_space[4414] = 8'h00;
reg_space[4415] = 8'h00;
reg_space[4416] = 8'h00;
reg_space[4417] = 8'h00;
reg_space[4418] = 8'h00;
reg_space[4419] = 8'h00;
reg_space[4420] = 8'h00;
reg_space[4421] = 8'h00;
reg_space[4422] = 8'h00;
reg_space[4423] = 8'h00;
reg_space[4424] = 8'h00;
reg_space[4425] = 8'h00;
reg_space[4426] = 8'h00;
reg_space[4427] = 8'h00;
reg_space[4428] = 8'h00;
reg_space[4429] = 8'h00;
reg_space[4430] = 8'h00;
reg_space[4431] = 8'h00;
reg_space[4432] = 8'h00;
reg_space[4433] = 8'h00;
reg_space[4434] = 8'h00;
reg_space[4435] = 8'h00;
reg_space[4436] = 8'h00;
reg_space[4437] = 8'h00;
reg_space[4438] = 8'h00;
reg_space[4439] = 8'h00;
reg_space[4440] = 8'h00;
reg_space[4441] = 8'h00;
reg_space[4442] = 8'h00;
reg_space[4443] = 8'h00;
reg_space[4444] = 8'h00;
reg_space[4445] = 8'h00;
reg_space[4446] = 8'h00;
reg_space[4447] = 8'h00;
reg_space[4448] = 8'h00;
reg_space[4449] = 8'h00;
reg_space[4450] = 8'h00;
reg_space[4451] = 8'h00;
reg_space[4452] = 8'h00;
reg_space[4453] = 8'h00;
reg_space[4454] = 8'h00;
reg_space[4455] = 8'h00;
reg_space[4456] = 8'h00;
reg_space[4457] = 8'h00;
reg_space[4458] = 8'h00;
reg_space[4459] = 8'h00;
reg_space[4460] = 8'h00;
reg_space[4461] = 8'h00;
reg_space[4462] = 8'h00;
reg_space[4463] = 8'h00;
reg_space[4464] = 8'h00;
reg_space[4465] = 8'h00;
reg_space[4466] = 8'h00;
reg_space[4467] = 8'h00;
reg_space[4468] = 8'h00;
reg_space[4469] = 8'h00;
reg_space[4470] = 8'h00;
reg_space[4471] = 8'h00;
reg_space[4472] = 8'h00;
reg_space[4473] = 8'h00;
reg_space[4474] = 8'h00;
reg_space[4475] = 8'h00;
reg_space[4476] = 8'h00;
reg_space[4477] = 8'h00;
reg_space[4478] = 8'h00;
reg_space[4479] = 8'h00;
reg_space[4480] = 8'h00;
reg_space[4481] = 8'h00;
reg_space[4482] = 8'h00;
reg_space[4483] = 8'h00;
reg_space[4484] = 8'h00;
reg_space[4485] = 8'h00;
reg_space[4486] = 8'h00;
reg_space[4487] = 8'h00;
reg_space[4488] = 8'h00;
reg_space[4489] = 8'h00;
reg_space[4490] = 8'h00;
reg_space[4491] = 8'h00;
reg_space[4492] = 8'h00;
reg_space[4493] = 8'h00;
reg_space[4494] = 8'h00;
reg_space[4495] = 8'h00;
reg_space[4496] = 8'h00;
reg_space[4497] = 8'h00;
reg_space[4498] = 8'h00;
reg_space[4499] = 8'h00;
reg_space[4500; = 8'h00;
reg_space[4501] = 8'h00;
reg_space[4502] = 8'h00;
reg_space[4503] = 8'h00;
reg_space[4504] = 8'h00;
reg_space[4505] = 8'h00;
reg_space[4506] = 8'h00;
reg_space[4507] = 8'h00;
reg_space[4508] = 8'h00;
reg_space[4509] = 8'h00;
reg_space[4510] = 8'h00;
reg_space[4511] = 8'h00;
reg_space[4512] = 8'h00;
reg_space[4513] = 8'h00;
reg_space[4514] = 8'h00;
reg_space[4515] = 8'h00;
reg_space[4516] = 8'h00;
reg_space[4517] = 8'h00;
reg_space[4518] = 8'h00;
reg_space[4519] = 8'h00;
reg_space[4520] = 8'h00;
reg_space[4521] = 8'h00;
reg_space[4522] = 8'h00;
reg_space[4523] = 8'h00;
reg_space[4524] = 8'h00;
reg_space[4525] = 8'h00;
reg_space[4526] = 8'h00;
reg_space[4527] = 8'h00;
reg_space[4528] = 8'h00;
reg_space[4529] = 8'h00;
reg_space[4530] = 8'h00;
reg_space[4531] = 8'h00;
reg_space[4532] = 8'h00;
reg_space[4533] = 8'h00;
reg_space[4534] = 8'h00;
reg_space[4535] = 8'h00;
reg_space[4536] = 8'h00;
reg_space[4537] = 8'h00;
reg_space[4538] = 8'h00;
reg_space[4539] = 8'h00;
reg_space[4540] = 8'h00;
reg_space[4541] = 8'h00;
reg_space[4542] = 8'h00;
reg_space[4543] = 8'h00;
reg_space[4544] = 8'h00;
reg_space[4545] = 8'h00;
reg_space[4546] = 8'h00;
reg_space[4547] = 8'h00;
reg_space[4548] = 8'h00;
reg_space[4549] = 8'h00;
reg_space[4550] = 8'h00;
reg_space[4551] = 8'h00;
reg_space[4552] = 8'h00;
reg_space[4553] = 8'h00;
reg_space[4554] = 8'h00;
reg_space[4555] = 8'h00;
reg_space[4556] = 8'h00;
reg_space[4557] = 8'h00;
reg_space[4558] = 8'h00;
reg_space[4559] = 8'h00;
reg_space[4560] = 8'h00;
reg_space[4561] = 8'h00;
reg_space[4562] = 8'h00;
reg_space[4563] = 8'h00;
reg_space[4564] = 8'h00;
reg_space[4565] = 8'h00;
reg_space[4566] = 8'h00;
reg_space[4567] = 8'h00;
reg_space[4568] = 8'h00;
reg_space[4569] = 8'h00;
reg_space[4570] = 8'h00;
reg_space[4571] = 8'h00;
reg_space[4572] = 8'h00;
reg_space[4573] = 8'h00;
reg_space[4574] = 8'h00;
reg_space[4575] = 8'h00;
reg_space[4576] = 8'h00;
reg_space[4577] = 8'h00;
reg_space[4578] = 8'h00;
reg_space[4579] = 8'h00;
reg_space[4580] = 8'h00;
reg_space[4581] = 8'h00;
reg_space[4582] = 8'h00;
reg_space[4583] = 8'h00;
reg_space[4584] = 8'h00;
reg_space[4585] = 8'h00;
reg_space[4586] = 8'h00;
reg_space[4587] = 8'h00;
reg_space[4588] = 8'h00;
reg_space[4589] = 8'h00;
reg_space[4590] = 8'h00;
reg_space[4591] = 8'h00;
reg_space[4592] = 8'h00;
reg_space[4593] = 8'h00;
reg_space[4594] = 8'h00;
reg_space[4595] = 8'h00;
reg_space[4596] = 8'h00;
reg_space[4597] = 8'h00;
reg_space[4598] = 8'h00;
reg_space[4599] = 8'h00;
reg_space[4600; = 8'h00;
reg_space[4601] = 8'h00;
reg_space[4602] = 8'h00;
reg_space[4603] = 8'h00;
reg_space[4604] = 8'h00;
reg_space[4605] = 8'h00;
reg_space[4606] = 8'h00;
reg_space[4607] = 8'h00;
reg_space[4608] = 8'h00;
reg_space[4609] = 8'h00;
reg_space[4610] = 8'h00;
reg_space[4611] = 8'h00;
reg_space[4612] = 8'h00;
reg_space[4613] = 8'h00;
reg_space[4614] = 8'h00;
reg_space[4615] = 8'h00;
reg_space[4616] = 8'h00;
reg_space[4617] = 8'h00;
reg_space[4618] = 8'h00;
reg_space[4619] = 8'h00;
reg_space[4620] = 8'h00;
reg_space[4621] = 8'h00;
reg_space[4622] = 8'h00;
reg_space[4623] = 8'h00;
reg_space[4624] = 8'h00;
reg_space[4625] = 8'h00;
reg_space[4626] = 8'h00;
reg_space[4627] = 8'h00;
reg_space[4628] = 8'h00;
reg_space[4629] = 8'h00;
reg_space[4630] = 8'h00;
reg_space[4631] = 8'h00;
reg_space[4632] = 8'h00;
reg_space[4633] = 8'h00;
reg_space[4634] = 8'h00;
reg_space[4635] = 8'h00;
reg_space[4636] = 8'h00;
reg_space[4637] = 8'h00;
reg_space[4638] = 8'h00;
reg_space[4639] = 8'h00;
reg_space[4640] = 8'h00;
reg_space[4641] = 8'h00;
reg_space[4642] = 8'h00;
reg_space[4643] = 8'h00;
reg_space[4644] = 8'h00;
reg_space[4645] = 8'h00;
reg_space[4646] = 8'h00;
reg_space[4647] = 8'h00;
reg_space[4648] = 8'h00;
reg_space[4649] = 8'h00;
reg_space[4650] = 8'h00;
reg_space[4651] = 8'h00;
reg_space[4652] = 8'h00;
reg_space[4653] = 8'h00;
reg_space[4654] = 8'h00;
reg_space[4655] = 8'h00;
reg_space[4656] = 8'h00;
reg_space[4657] = 8'h00;
reg_space[4658] = 8'h00;
reg_space[4659] = 8'h00;
reg_space[4660] = 8'h00;
reg_space[4661] = 8'h00;
reg_space[4662] = 8'h00;
reg_space[4663] = 8'h00;
reg_space[4664] = 8'h00;
reg_space[4665] = 8'h00;
reg_space[4666] = 8'h00;
reg_space[4667] = 8'h00;
reg_space[4668] = 8'h00;
reg_space[4669] = 8'h00;
reg_space[4670] = 8'h00;
reg_space[4671] = 8'h00;
reg_space[4672] = 8'h00;
reg_space[4673] = 8'h00;
reg_space[4674] = 8'h00;
reg_space[4675] = 8'h00;
reg_space[4676] = 8'h00;
reg_space[4677] = 8'h00;
reg_space[4678] = 8'h00;
reg_space[4679] = 8'h00;
reg_space[4680] = 8'h00;
reg_space[4681] = 8'h00;
reg_space[4682] = 8'h00;
reg_space[4683] = 8'h00;
reg_space[4684] = 8'h00;
reg_space[4685] = 8'h00;
reg_space[4686] = 8'h00;
reg_space[4687] = 8'h00;
reg_space[4688] = 8'h00;
reg_space[4689] = 8'h00;
reg_space[4690] = 8'h00;
reg_space[4691] = 8'h00;
reg_space[4692] = 8'h00;
reg_space[4693] = 8'h00;
reg_space[4694] = 8'h00;
reg_space[4695] = 8'h00;
reg_space[4696] = 8'h00;
reg_space[4697] = 8'h00;
reg_space[4698] = 8'h00;
reg_space[4699] = 8'h00;
reg_space[4700; = 8'h00;
reg_space[4701] = 8'h00;
reg_space[4702] = 8'h00;
reg_space[4703] = 8'h00;
reg_space[4704] = 8'h00;
reg_space[4705] = 8'h00;
reg_space[4706] = 8'h00;
reg_space[4707] = 8'h00;
reg_space[4708] = 8'h00;
reg_space[4709] = 8'h00;
reg_space[4710] = 8'h00;
reg_space[4711] = 8'h00;
reg_space[4712] = 8'h00;
reg_space[4713] = 8'h00;
reg_space[4714] = 8'h00;
reg_space[4715] = 8'h00;
reg_space[4716] = 8'h00;
reg_space[4717] = 8'h00;
reg_space[4718] = 8'h00;
reg_space[4719] = 8'h00;
reg_space[4720] = 8'h00;
reg_space[4721] = 8'h00;
reg_space[4722] = 8'h00;
reg_space[4723] = 8'h00;
reg_space[4724] = 8'h00;
reg_space[4725] = 8'h00;
reg_space[4726] = 8'h00;
reg_space[4727] = 8'h00;
reg_space[4728] = 8'h00;
reg_space[4729] = 8'h00;
reg_space[4730] = 8'h00;
reg_space[4731] = 8'h00;
reg_space[4732] = 8'h00;
reg_space[4733] = 8'h00;
reg_space[4734] = 8'h00;
reg_space[4735] = 8'h00;
reg_space[4736] = 8'h00;
reg_space[4737] = 8'h00;
reg_space[4738] = 8'h00;
reg_space[4739] = 8'h00;
reg_space[4740] = 8'h00;
reg_space[4741] = 8'h00;
reg_space[4742] = 8'h00;
reg_space[4743] = 8'h00;
reg_space[4744] = 8'h00;
reg_space[4745] = 8'h00;
reg_space[4746] = 8'h00;
reg_space[4747] = 8'h00;
reg_space[4748] = 8'h00;
reg_space[4749] = 8'h00;
reg_space[4750] = 8'h00;
reg_space[4751] = 8'h00;
reg_space[4752] = 8'h00;
reg_space[4753] = 8'h00;
reg_space[4754] = 8'h00;
reg_space[4755] = 8'h00;
reg_space[4756] = 8'h00;
reg_space[4757] = 8'h00;
reg_space[4758] = 8'h00;
reg_space[4759] = 8'h00;
reg_space[4760] = 8'h00;
reg_space[4761] = 8'h00;
reg_space[4762] = 8'h00;
reg_space[4763] = 8'h00;
reg_space[4764] = 8'h00;
reg_space[4765] = 8'h00;
reg_space[4766] = 8'h00;
reg_space[4767] = 8'h00;
reg_space[4768] = 8'h00;
reg_space[4769] = 8'h00;
reg_space[4770] = 8'h00;
reg_space[4771] = 8'h00;
reg_space[4772] = 8'h00;
reg_space[4773] = 8'h00;
reg_space[4774] = 8'h00;
reg_space[4775] = 8'h00;
reg_space[4776] = 8'h00;
reg_space[4777] = 8'h00;
reg_space[4778] = 8'h00;
reg_space[4779] = 8'h00;
reg_space[4780] = 8'h00;
reg_space[4781] = 8'h00;
reg_space[4782] = 8'h00;
reg_space[4783] = 8'h00;
reg_space[4784] = 8'h00;
reg_space[4785] = 8'h00;
reg_space[4786] = 8'h00;
reg_space[4787] = 8'h00;
reg_space[4788] = 8'h00;
reg_space[4789] = 8'h00;
reg_space[4790] = 8'h00;
reg_space[4791] = 8'h00;
reg_space[4792] = 8'h00;
reg_space[4793] = 8'h00;
reg_space[4794] = 8'h00;
reg_space[4795] = 8'h00;
reg_space[4796] = 8'h00;
reg_space[4797] = 8'h00;
reg_space[4798] = 8'h00;
reg_space[4799] = 8'h00;
reg_space[4800; = 8'h00;
reg_space[4801] = 8'h00;
reg_space[4802] = 8'h00;
reg_space[4803] = 8'h00;
reg_space[4804] = 8'h00;
reg_space[4805] = 8'h00;
reg_space[4806] = 8'h00;
reg_space[4807] = 8'h00;
reg_space[4808] = 8'h00;
reg_space[4809] = 8'h00;
reg_space[4810] = 8'h00;
reg_space[4811] = 8'h00;
reg_space[4812] = 8'h00;
reg_space[4813] = 8'h00;
reg_space[4814] = 8'h00;
reg_space[4815] = 8'h00;
reg_space[4816] = 8'h00;
reg_space[4817] = 8'h00;
reg_space[4818] = 8'h00;
reg_space[4819] = 8'h00;
reg_space[4820] = 8'h00;
reg_space[4821] = 8'h00;
reg_space[4822] = 8'h00;
reg_space[4823] = 8'h00;
reg_space[4824] = 8'h00;
reg_space[4825] = 8'h00;
reg_space[4826] = 8'h00;
reg_space[4827] = 8'h00;
reg_space[4828] = 8'h00;
reg_space[4829] = 8'h00;
reg_space[4830] = 8'h00;
reg_space[4831] = 8'h00;
reg_space[4832] = 8'h00;
reg_space[4833] = 8'h00;
reg_space[4834] = 8'h00;
reg_space[4835] = 8'h00;
reg_space[4836] = 8'h00;
reg_space[4837] = 8'h00;
reg_space[4838] = 8'h00;
reg_space[4839] = 8'h00;
reg_space[4840] = 8'h00;
reg_space[4841] = 8'h00;
reg_space[4842] = 8'h00;
reg_space[4843] = 8'h00;
reg_space[4844] = 8'h00;
reg_space[4845] = 8'h00;
reg_space[4846] = 8'h00;
reg_space[4847] = 8'h00;
reg_space[4848] = 8'h00;
reg_space[4849] = 8'h00;
reg_space[4850] = 8'h00;
reg_space[4851] = 8'h00;
reg_space[4852] = 8'h00;
reg_space[4853] = 8'h00;
reg_space[4854] = 8'h00;
reg_space[4855] = 8'h00;
reg_space[4856] = 8'h00;
reg_space[4857] = 8'h00;
reg_space[4858] = 8'h00;
reg_space[4859] = 8'h00;
reg_space[4860] = 8'h00;
reg_space[4861] = 8'h00;
reg_space[4862] = 8'h00;
reg_space[4863] = 8'h00;
reg_space[4864] = 8'h00;
reg_space[4865] = 8'h00;
reg_space[4866] = 8'h00;
reg_space[4867] = 8'h00;
reg_space[4868] = 8'h00;
reg_space[4869] = 8'h00;
reg_space[4870] = 8'h00;
reg_space[4871] = 8'h00;
reg_space[4872] = 8'h00;
reg_space[4873] = 8'h00;
reg_space[4874] = 8'h00;
reg_space[4875] = 8'h00;
reg_space[4876] = 8'h00;
reg_space[4877] = 8'h00;
reg_space[4878] = 8'h00;
reg_space[4879] = 8'h00;
reg_space[4880] = 8'h00;
reg_space[4881] = 8'h00;
reg_space[4882] = 8'h00;
reg_space[4883] = 8'h00;
reg_space[4884] = 8'h00;
reg_space[4885] = 8'h00;
reg_space[4886] = 8'h00;
reg_space[4887] = 8'h00;
reg_space[4888] = 8'h00;
reg_space[4889] = 8'h00;
reg_space[4890] = 8'h00;
reg_space[4891] = 8'h00;
reg_space[4892] = 8'h00;
reg_space[4893] = 8'h00;
reg_space[4894] = 8'h00;
reg_space[4895] = 8'h00;
reg_space[4896] = 8'h00;
reg_space[4897] = 8'h00;
reg_space[4898] = 8'h00;
reg_space[4899] = 8'h00;
reg_space[4900; = 8'h00;
reg_space[4901] = 8'h00;
reg_space[4902] = 8'h00;
reg_space[4903] = 8'h00;
reg_space[4904] = 8'h00;
reg_space[4905] = 8'h00;
reg_space[4906] = 8'h00;
reg_space[4907] = 8'h00;
reg_space[4908] = 8'h00;
reg_space[4909] = 8'h00;
reg_space[4910] = 8'h00;
reg_space[4911] = 8'h00;
reg_space[4912] = 8'h00;
reg_space[4913] = 8'h00;
reg_space[4914] = 8'h00;
reg_space[4915] = 8'h00;
reg_space[4916] = 8'h00;
reg_space[4917] = 8'h00;
reg_space[4918] = 8'h00;
reg_space[4919] = 8'h00;
reg_space[4920] = 8'h00;
reg_space[4921] = 8'h00;
reg_space[4922] = 8'h00;
reg_space[4923] = 8'h00;
reg_space[4924] = 8'h00;
reg_space[4925] = 8'h00;
reg_space[4926] = 8'h00;
reg_space[4927] = 8'h00;
reg_space[4928] = 8'h00;
reg_space[4929] = 8'h00;
reg_space[4930] = 8'h00;
reg_space[4931] = 8'h00;
reg_space[4932] = 8'h00;
reg_space[4933] = 8'h00;
reg_space[4934] = 8'h00;
reg_space[4935] = 8'h00;
reg_space[4936] = 8'h00;
reg_space[4937] = 8'h00;
reg_space[4938] = 8'h00;
reg_space[4939] = 8'h00;
reg_space[4940] = 8'h00;
reg_space[4941] = 8'h00;
reg_space[4942] = 8'h00;
reg_space[4943] = 8'h00;
reg_space[4944] = 8'h00;
reg_space[4945] = 8'h00;
reg_space[4946] = 8'h00;
reg_space[4947] = 8'h00;
reg_space[4948] = 8'h00;
reg_space[4949] = 8'h00;
reg_space[4950] = 8'h00;
reg_space[4951] = 8'h00;
reg_space[4952] = 8'h00;
reg_space[4953] = 8'h00;
reg_space[4954] = 8'h00;
reg_space[4955] = 8'h00;
reg_space[4956] = 8'h00;
reg_space[4957] = 8'h00;
reg_space[4958] = 8'h00;
reg_space[4959] = 8'h00;
reg_space[4960] = 8'h00;
reg_space[4961] = 8'h00;
reg_space[4962] = 8'h00;
reg_space[4963] = 8'h00;
reg_space[4964] = 8'h00;
reg_space[4965] = 8'h00;
reg_space[4966] = 8'h00;
reg_space[4967] = 8'h00;
reg_space[4968] = 8'h00;
reg_space[4969] = 8'h00;
reg_space[4970] = 8'h00;
reg_space[4971] = 8'h00;
reg_space[4972] = 8'h00;
reg_space[4973] = 8'h00;
reg_space[4974] = 8'h00;
reg_space[4975] = 8'h00;
reg_space[4976] = 8'h00;
reg_space[4977] = 8'h00;
reg_space[4978] = 8'h00;
reg_space[4979] = 8'h00;
reg_space[4980] = 8'h00;
reg_space[4981] = 8'h00;
reg_space[4982] = 8'h00;
reg_space[4983] = 8'h00;
reg_space[4984] = 8'h00;
reg_space[4985] = 8'h00;
reg_space[4986] = 8'h00;
reg_space[4987] = 8'h00;
reg_space[4988] = 8'h00;
reg_space[4989] = 8'h00;
reg_space[4990] = 8'h00;
reg_space[4991] = 8'h00;
reg_space[4992] = 8'h00;
reg_space[4993] = 8'h00;
reg_space[4994] = 8'h00;
reg_space[4995] = 8'h00;
reg_space[4996] = 8'h00;
reg_space[4997] = 8'h00;
reg_space[4998] = 8'h00;
reg_space[4999] = 8'h00;
reg_space[500;0] = 8'h00;
reg_space[500;1] = 8'h00;
reg_space[500;2] = 8'h00;
reg_space[500;3] = 8'h00;
reg_space[500;4] = 8'h00;
reg_space[500;5] = 8'h00;
reg_space[500;6] = 8'h00;
reg_space[500;7] = 8'h00;
reg_space[500;8] = 8'h00;
reg_space[500;9] = 8'h00;
reg_space[5010] = 8'h00;
reg_space[5011] = 8'h00;
reg_space[5012] = 8'h00;
reg_space[5013] = 8'h00;
reg_space[5014] = 8'h00;
reg_space[5015] = 8'h00;
reg_space[5016] = 8'h00;
reg_space[5017] = 8'h00;
reg_space[5018] = 8'h00;
reg_space[5019] = 8'h00;
reg_space[5020] = 8'h00;
reg_space[5021] = 8'h00;
reg_space[5022] = 8'h00;
reg_space[5023] = 8'h00;
reg_space[5024] = 8'h00;
reg_space[5025] = 8'h00;
reg_space[5026] = 8'h00;
reg_space[5027] = 8'h00;
reg_space[5028] = 8'h00;
reg_space[5029] = 8'h00;
reg_space[5030] = 8'h00;
reg_space[5031] = 8'h00;
reg_space[5032] = 8'h00;
reg_space[5033] = 8'h00;
reg_space[5034] = 8'h00;
reg_space[5035] = 8'h00;
reg_space[5036] = 8'h00;
reg_space[5037] = 8'h00;
reg_space[5038] = 8'h00;
reg_space[5039] = 8'h00;
reg_space[5040] = 8'h00;
reg_space[5041] = 8'h00;
reg_space[5042] = 8'h00;
reg_space[5043] = 8'h00;
reg_space[5044] = 8'h00;
reg_space[5045] = 8'h00;
reg_space[5046] = 8'h00;
reg_space[5047] = 8'h00;
reg_space[5048] = 8'h00;
reg_space[5049] = 8'h00;
reg_space[5050] = 8'h00;
reg_space[5051] = 8'h00;
reg_space[5052] = 8'h00;
reg_space[5053] = 8'h00;
reg_space[5054] = 8'h00;
reg_space[5055] = 8'h00;
reg_space[5056] = 8'h00;
reg_space[5057] = 8'h00;
reg_space[5058] = 8'h00;
reg_space[5059] = 8'h00;
reg_space[5060] = 8'h00;
reg_space[5061] = 8'h00;
reg_space[5062] = 8'h00;
reg_space[5063] = 8'h00;
reg_space[5064] = 8'h00;
reg_space[5065] = 8'h00;
reg_space[5066] = 8'h00;
reg_space[5067] = 8'h00;
reg_space[5068] = 8'h00;
reg_space[5069] = 8'h00;
reg_space[5070] = 8'h00;
reg_space[5071] = 8'h00;
reg_space[5072] = 8'h00;
reg_space[5073] = 8'h00;
reg_space[5074] = 8'h00;
reg_space[5075] = 8'h00;
reg_space[5076] = 8'h00;
reg_space[5077] = 8'h00;
reg_space[5078] = 8'h00;
reg_space[5079] = 8'h00;
reg_space[5080] = 8'h00;
reg_space[5081] = 8'h00;
reg_space[5082] = 8'h00;
reg_space[5083] = 8'h00;
reg_space[5084] = 8'h00;
reg_space[5085] = 8'h00;
reg_space[5086] = 8'h00;
reg_space[5087] = 8'h00;
reg_space[5088] = 8'h00;
reg_space[5089] = 8'h00;
reg_space[5090] = 8'h00;
reg_space[5091] = 8'h00;
reg_space[5092] = 8'h00;
reg_space[5093] = 8'h00;
reg_space[5094] = 8'h00;
reg_space[5095] = 8'h00;
reg_space[5096] = 8'h00;
reg_space[5097] = 8'h00;
reg_space[5098] = 8'h00;
reg_space[5099] = 8'h00;
reg_space[5100; = 8'h00;
reg_space[5101] = 8'h00;
reg_space[5102] = 8'h00;
reg_space[5103] = 8'h00;
reg_space[5104] = 8'h00;
reg_space[5105] = 8'h00;
reg_space[5106] = 8'h00;
reg_space[5107] = 8'h00;
reg_space[5108] = 8'h00;
reg_space[5109] = 8'h00;
reg_space[5110] = 8'h00;
reg_space[5111] = 8'h00;
reg_space[5112] = 8'h00;
reg_space[5113] = 8'h00;
reg_space[5114] = 8'h00;
reg_space[5115] = 8'h00;
reg_space[5116] = 8'h00;
reg_space[5117] = 8'h00;
reg_space[5118] = 8'h00;
reg_space[5119] = 8'h00;
reg_space[5120] = 8'h00;
reg_space[5121] = 8'h00;
reg_space[5122] = 8'h00;
reg_space[5123] = 8'h00;
reg_space[5124] = 8'h00;
reg_space[5125] = 8'h00;
reg_space[5126] = 8'h00;
reg_space[5127] = 8'h00;
reg_space[5128] = 8'h00;
reg_space[5129] = 8'h00;
reg_space[5130] = 8'h00;
reg_space[5131] = 8'h00;
reg_space[5132] = 8'h00;
reg_space[5133] = 8'h00;
reg_space[5134] = 8'h00;
reg_space[5135] = 8'h00;
reg_space[5136] = 8'h00;
reg_space[5137] = 8'h00;
reg_space[5138] = 8'h00;
reg_space[5139] = 8'h00;
reg_space[5140] = 8'h00;
reg_space[5141] = 8'h00;
reg_space[5142] = 8'h00;
reg_space[5143] = 8'h00;
reg_space[5144] = 8'h00;
reg_space[5145] = 8'h00;
reg_space[5146] = 8'h00;
reg_space[5147] = 8'h00;
reg_space[5148] = 8'h00;
reg_space[5149] = 8'h00;
reg_space[5150] = 8'h00;
reg_space[5151] = 8'h00;
reg_space[5152] = 8'h00;
reg_space[5153] = 8'h00;
reg_space[5154] = 8'h00;
reg_space[5155] = 8'h00;
reg_space[5156] = 8'h00;
reg_space[5157] = 8'h00;
reg_space[5158] = 8'h00;
reg_space[5159] = 8'h00;
reg_space[5160] = 8'h00;
reg_space[5161] = 8'h00;
reg_space[5162] = 8'h00;
reg_space[5163] = 8'h00;
reg_space[5164] = 8'h00;
reg_space[5165] = 8'h00;
reg_space[5166] = 8'h00;
reg_space[5167] = 8'h00;
reg_space[5168] = 8'h00;
reg_space[5169] = 8'h00;
reg_space[5170] = 8'h00;
reg_space[5171] = 8'h00;
reg_space[5172] = 8'h00;
reg_space[5173] = 8'h00;
reg_space[5174] = 8'h00;
reg_space[5175] = 8'h00;
reg_space[5176] = 8'h00;
reg_space[5177] = 8'h00;
reg_space[5178] = 8'h00;
reg_space[5179] = 8'h00;
reg_space[5180] = 8'h00;
reg_space[5181] = 8'h00;
reg_space[5182] = 8'h00;
reg_space[5183] = 8'h00;
reg_space[5184] = 8'h00;
reg_space[5185] = 8'h00;
reg_space[5186] = 8'h00;
reg_space[5187] = 8'h00;
reg_space[5188] = 8'h00;
reg_space[5189] = 8'h00;
reg_space[5190] = 8'h00;
reg_space[5191] = 8'h00;
reg_space[5192] = 8'h00;
reg_space[5193] = 8'h00;
reg_space[5194] = 8'h00;
reg_space[5195] = 8'h00;
reg_space[5196] = 8'h00;
reg_space[5197] = 8'h00;
reg_space[5198] = 8'h00;
reg_space[5199] = 8'h00;
reg_space[5200; = 8'h00;
reg_space[5201] = 8'h00;
reg_space[5202] = 8'h00;
reg_space[5203] = 8'h00;
reg_space[5204] = 8'h00;
reg_space[5205] = 8'h00;
reg_space[5206] = 8'h00;
reg_space[5207] = 8'h00;
reg_space[5208] = 8'h00;
reg_space[5209] = 8'h00;
reg_space[5210] = 8'h00;
reg_space[5211] = 8'h00;
reg_space[5212] = 8'h00;
reg_space[5213] = 8'h00;
reg_space[5214] = 8'h00;
reg_space[5215] = 8'h00;
reg_space[5216] = 8'h00;
reg_space[5217] = 8'h00;
reg_space[5218] = 8'h00;
reg_space[5219] = 8'h00;
reg_space[5220] = 8'h00;
reg_space[5221] = 8'h00;
reg_space[5222] = 8'h00;
reg_space[5223] = 8'h00;
reg_space[5224] = 8'h00;
reg_space[5225] = 8'h00;
reg_space[5226] = 8'h00;
reg_space[5227] = 8'h00;
reg_space[5228] = 8'h00;
reg_space[5229] = 8'h00;
reg_space[5230] = 8'h00;
reg_space[5231] = 8'h00;
reg_space[5232] = 8'h00;
reg_space[5233] = 8'h00;
reg_space[5234] = 8'h00;
reg_space[5235] = 8'h00;
reg_space[5236] = 8'h00;
reg_space[5237] = 8'h00;
reg_space[5238] = 8'h00;
reg_space[5239] = 8'h00;
reg_space[5240] = 8'h00;
reg_space[5241] = 8'h00;
reg_space[5242] = 8'h00;
reg_space[5243] = 8'h00;
reg_space[5244] = 8'h00;
reg_space[5245] = 8'h00;
reg_space[5246] = 8'h00;
reg_space[5247] = 8'h00;
reg_space[5248] = 8'h00;
reg_space[5249] = 8'h00;
reg_space[5250] = 8'h00;
reg_space[5251] = 8'h00;
reg_space[5252] = 8'h00;
reg_space[5253] = 8'h00;
reg_space[5254] = 8'h00;
reg_space[5255] = 8'h00;
reg_space[5256] = 8'h00;
reg_space[5257] = 8'h00;
reg_space[5258] = 8'h00;
reg_space[5259] = 8'h00;
reg_space[5260] = 8'h00;
reg_space[5261] = 8'h00;
reg_space[5262] = 8'h00;
reg_space[5263] = 8'h00;
reg_space[5264] = 8'h00;
reg_space[5265] = 8'h00;
reg_space[5266] = 8'h00;
reg_space[5267] = 8'h00;
reg_space[5268] = 8'h00;
reg_space[5269] = 8'h00;
reg_space[5270] = 8'h00;
reg_space[5271] = 8'h00;
reg_space[5272] = 8'h00;
reg_space[5273] = 8'h00;
reg_space[5274] = 8'h00;
reg_space[5275] = 8'h00;
reg_space[5276] = 8'h00;
reg_space[5277] = 8'h00;
reg_space[5278] = 8'h00;
reg_space[5279] = 8'h00;
reg_space[5280] = 8'h00;
reg_space[5281] = 8'h00;
reg_space[5282] = 8'h00;
reg_space[5283] = 8'h00;
reg_space[5284] = 8'h00;
reg_space[5285] = 8'h00;
reg_space[5286] = 8'h00;
reg_space[5287] = 8'h00;
reg_space[5288] = 8'h00;
reg_space[5289] = 8'h00;
reg_space[5290] = 8'h00;
reg_space[5291] = 8'h00;
reg_space[5292] = 8'h00;
reg_space[5293] = 8'h00;
reg_space[5294] = 8'h00;
reg_space[5295] = 8'h00;
reg_space[5296] = 8'h00;
reg_space[5297] = 8'h00;
reg_space[5298] = 8'h00;
reg_space[5299] = 8'h00;
reg_space[5300; = 8'h00;
reg_space[5301] = 8'h00;
reg_space[5302] = 8'h00;
reg_space[5303] = 8'h00;
reg_space[5304] = 8'h00;
reg_space[5305] = 8'h00;
reg_space[5306] = 8'h00;
reg_space[5307] = 8'h00;
reg_space[5308] = 8'h00;
reg_space[5309] = 8'h00;
reg_space[5310] = 8'h00;
reg_space[5311] = 8'h00;
reg_space[5312] = 8'h00;
reg_space[5313] = 8'h00;
reg_space[5314] = 8'h00;
reg_space[5315] = 8'h00;
reg_space[5316] = 8'h00;
reg_space[5317] = 8'h00;
reg_space[5318] = 8'h00;
reg_space[5319] = 8'h00;
reg_space[5320] = 8'h00;
reg_space[5321] = 8'h00;
reg_space[5322] = 8'h00;
reg_space[5323] = 8'h00;
reg_space[5324] = 8'h00;
reg_space[5325] = 8'h00;
reg_space[5326] = 8'h00;
reg_space[5327] = 8'h00;
reg_space[5328] = 8'h00;
reg_space[5329] = 8'h00;
reg_space[5330] = 8'h00;
reg_space[5331] = 8'h00;
reg_space[5332] = 8'h00;
reg_space[5333] = 8'h00;
reg_space[5334] = 8'h00;
reg_space[5335] = 8'h00;
reg_space[5336] = 8'h00;
reg_space[5337] = 8'h00;
reg_space[5338] = 8'h00;
reg_space[5339] = 8'h00;
reg_space[5340] = 8'h00;
reg_space[5341] = 8'h00;
reg_space[5342] = 8'h00;
reg_space[5343] = 8'h00;
reg_space[5344] = 8'h00;
reg_space[5345] = 8'h00;
reg_space[5346] = 8'h00;
reg_space[5347] = 8'h00;
reg_space[5348] = 8'h00;
reg_space[5349] = 8'h00;
reg_space[5350] = 8'h00;
reg_space[5351] = 8'h00;
reg_space[5352] = 8'h00;
reg_space[5353] = 8'h00;
reg_space[5354] = 8'h00;
reg_space[5355] = 8'h00;
reg_space[5356] = 8'h00;
reg_space[5357] = 8'h00;
reg_space[5358] = 8'h00;
reg_space[5359] = 8'h00;
reg_space[5360] = 8'h00;
reg_space[5361] = 8'h00;
reg_space[5362] = 8'h00;
reg_space[5363] = 8'h00;
reg_space[5364] = 8'h00;
reg_space[5365] = 8'h00;
reg_space[5366] = 8'h00;
reg_space[5367] = 8'h00;
reg_space[5368] = 8'h00;
reg_space[5369] = 8'h00;
reg_space[5370] = 8'h00;
reg_space[5371] = 8'h00;
reg_space[5372] = 8'h00;
reg_space[5373] = 8'h00;
reg_space[5374] = 8'h00;
reg_space[5375] = 8'h00;
reg_space[5376] = 8'h00;
reg_space[5377] = 8'h00;
reg_space[5378] = 8'h00;
reg_space[5379] = 8'h00;
reg_space[5380] = 8'h00;
reg_space[5381] = 8'h00;
reg_space[5382] = 8'h00;
reg_space[5383] = 8'h00;
reg_space[5384] = 8'h00;
reg_space[5385] = 8'h00;
reg_space[5386] = 8'h00;
reg_space[5387] = 8'h00;
reg_space[5388] = 8'h00;
reg_space[5389] = 8'h00;
reg_space[5390] = 8'h00;
reg_space[5391] = 8'h00;
reg_space[5392] = 8'h00;
reg_space[5393] = 8'h00;
reg_space[5394] = 8'h00;
reg_space[5395] = 8'h00;
reg_space[5396] = 8'h00;
reg_space[5397] = 8'h00;
reg_space[5398] = 8'h00;
reg_space[5399] = 8'h00;
reg_space[5400; = 8'h00;
reg_space[5401] = 8'h00;
reg_space[5402] = 8'h00;
reg_space[5403] = 8'h00;
reg_space[5404] = 8'h00;
reg_space[5405] = 8'h00;
reg_space[5406] = 8'h00;
reg_space[5407] = 8'h00;
reg_space[5408] = 8'h00;
reg_space[5409] = 8'h00;
reg_space[5410] = 8'h00;
reg_space[5411] = 8'h00;
reg_space[5412] = 8'h00;
reg_space[5413] = 8'h00;
reg_space[5414] = 8'h00;
reg_space[5415] = 8'h00;
reg_space[5416] = 8'h00;
reg_space[5417] = 8'h00;
reg_space[5418] = 8'h00;
reg_space[5419] = 8'h00;
reg_space[5420] = 8'h00;
reg_space[5421] = 8'h00;
reg_space[5422] = 8'h00;
reg_space[5423] = 8'h00;
reg_space[5424] = 8'h00;
reg_space[5425] = 8'h00;
reg_space[5426] = 8'h00;
reg_space[5427] = 8'h00;
reg_space[5428] = 8'h00;
reg_space[5429] = 8'h00;
reg_space[5430] = 8'h00;
reg_space[5431] = 8'h00;
reg_space[5432] = 8'h00;
reg_space[5433] = 8'h00;
reg_space[5434] = 8'h00;
reg_space[5435] = 8'h00;
reg_space[5436] = 8'h00;
reg_space[5437] = 8'h00;
reg_space[5438] = 8'h00;
reg_space[5439] = 8'h00;
reg_space[5440] = 8'h00;
reg_space[5441] = 8'h00;
reg_space[5442] = 8'h00;
reg_space[5443] = 8'h00;
reg_space[5444] = 8'h00;
reg_space[5445] = 8'h00;
reg_space[5446] = 8'h00;
reg_space[5447] = 8'h00;
reg_space[5448] = 8'h00;
reg_space[5449] = 8'h00;
reg_space[5450] = 8'h00;
reg_space[5451] = 8'h00;
reg_space[5452] = 8'h00;
reg_space[5453] = 8'h00;
reg_space[5454] = 8'h00;
reg_space[5455] = 8'h00;
reg_space[5456] = 8'h00;
reg_space[5457] = 8'h00;
reg_space[5458] = 8'h00;
reg_space[5459] = 8'h00;
reg_space[5460] = 8'h00;
reg_space[5461] = 8'h00;
reg_space[5462] = 8'h00;
reg_space[5463] = 8'h00;
reg_space[5464] = 8'h00;
reg_space[5465] = 8'h00;
reg_space[5466] = 8'h00;
reg_space[5467] = 8'h00;
reg_space[5468] = 8'h00;
reg_space[5469] = 8'h00;
reg_space[5470] = 8'h00;
reg_space[5471] = 8'h00;
reg_space[5472] = 8'h00;
reg_space[5473] = 8'h00;
reg_space[5474] = 8'h00;
reg_space[5475] = 8'h00;
reg_space[5476] = 8'h00;
reg_space[5477] = 8'h00;
reg_space[5478] = 8'h00;
reg_space[5479] = 8'h00;
reg_space[5480] = 8'h00;
reg_space[5481] = 8'h00;
reg_space[5482] = 8'h00;
reg_space[5483] = 8'h00;
reg_space[5484] = 8'h00;
reg_space[5485] = 8'h00;
reg_space[5486] = 8'h00;
reg_space[5487] = 8'h00;
reg_space[5488] = 8'h00;
reg_space[5489] = 8'h00;
reg_space[5490] = 8'h00;
reg_space[5491] = 8'h00;
reg_space[5492] = 8'h00;
reg_space[5493] = 8'h00;
reg_space[5494] = 8'h00;
reg_space[5495] = 8'h00;
reg_space[5496] = 8'h00;
reg_space[5497] = 8'h00;
reg_space[5498] = 8'h00;
reg_space[5499] = 8'h00;
reg_space[5500; = 8'h00;
reg_space[5501] = 8'h00;
reg_space[5502] = 8'h00;
reg_space[5503] = 8'h00;
reg_space[5504] = 8'h00;
reg_space[5505] = 8'h00;
reg_space[5506] = 8'h00;
reg_space[5507] = 8'h00;
reg_space[5508] = 8'h00;
reg_space[5509] = 8'h00;
reg_space[5510] = 8'h00;
reg_space[5511] = 8'h00;
reg_space[5512] = 8'h00;
reg_space[5513] = 8'h00;
reg_space[5514] = 8'h00;
reg_space[5515] = 8'h00;
reg_space[5516] = 8'h00;
reg_space[5517] = 8'h00;
reg_space[5518] = 8'h00;
reg_space[5519] = 8'h00;
reg_space[5520] = 8'h00;
reg_space[5521] = 8'h00;
reg_space[5522] = 8'h00;
reg_space[5523] = 8'h00;
reg_space[5524] = 8'h00;
reg_space[5525] = 8'h00;
reg_space[5526] = 8'h00;
reg_space[5527] = 8'h00;
reg_space[5528] = 8'h00;
reg_space[5529] = 8'h00;
reg_space[5530] = 8'h00;
reg_space[5531] = 8'h00;
reg_space[5532] = 8'h00;
reg_space[5533] = 8'h00;
reg_space[5534] = 8'h00;
reg_space[5535] = 8'h00;
reg_space[5536] = 8'h00;
reg_space[5537] = 8'h00;
reg_space[5538] = 8'h00;
reg_space[5539] = 8'h00;
reg_space[5540] = 8'h00;
reg_space[5541] = 8'h00;
reg_space[5542] = 8'h00;
reg_space[5543] = 8'h00;
reg_space[5544] = 8'h00;
reg_space[5545] = 8'h00;
reg_space[5546] = 8'h00;
reg_space[5547] = 8'h00;
reg_space[5548] = 8'h00;
reg_space[5549] = 8'h00;
reg_space[5550] = 8'h00;
reg_space[5551] = 8'h00;
reg_space[5552] = 8'h00;
reg_space[5553] = 8'h00;
reg_space[5554] = 8'h00;
reg_space[5555] = 8'h00;
reg_space[5556] = 8'h00;
reg_space[5557] = 8'h00;
reg_space[5558] = 8'h00;
reg_space[5559] = 8'h00;
reg_space[5560] = 8'h00;
reg_space[5561] = 8'h00;
reg_space[5562] = 8'h00;
reg_space[5563] = 8'h00;
reg_space[5564] = 8'h00;
reg_space[5565] = 8'h00;
reg_space[5566] = 8'h00;
reg_space[5567] = 8'h00;
reg_space[5568] = 8'h00;
reg_space[5569] = 8'h00;
reg_space[5570] = 8'h00;
reg_space[5571] = 8'h00;
reg_space[5572] = 8'h00;
reg_space[5573] = 8'h00;
reg_space[5574] = 8'h00;
reg_space[5575] = 8'h00;
reg_space[5576] = 8'h00;
reg_space[5577] = 8'h00;
reg_space[5578] = 8'h00;
reg_space[5579] = 8'h00;
reg_space[5580] = 8'h00;
reg_space[5581] = 8'h00;
reg_space[5582] = 8'h00;
reg_space[5583] = 8'h00;
reg_space[5584] = 8'h00;
reg_space[5585] = 8'h00;
reg_space[5586] = 8'h00;
reg_space[5587] = 8'h00;
reg_space[5588] = 8'h00;
reg_space[5589] = 8'h00;
reg_space[5590] = 8'h00;
reg_space[5591] = 8'h00;
reg_space[5592] = 8'h00;
reg_space[5593] = 8'h00;
reg_space[5594] = 8'h00;
reg_space[5595] = 8'h00;
reg_space[5596] = 8'h00;
reg_space[5597] = 8'h00;
reg_space[5598] = 8'h00;
reg_space[5599] = 8'h00;
reg_space[5600; = 8'h00;
reg_space[5601] = 8'h00;
reg_space[5602] = 8'h00;
reg_space[5603] = 8'h00;
reg_space[5604] = 8'h00;
reg_space[5605] = 8'h00;
reg_space[5606] = 8'h00;
reg_space[5607] = 8'h00;
reg_space[5608] = 8'h00;
reg_space[5609] = 8'h00;
reg_space[5610] = 8'h00;
reg_space[5611] = 8'h00;
reg_space[5612] = 8'h00;
reg_space[5613] = 8'h00;
reg_space[5614] = 8'h00;
reg_space[5615] = 8'h00;
reg_space[5616] = 8'h00;
reg_space[5617] = 8'h00;
reg_space[5618] = 8'h00;
reg_space[5619] = 8'h00;
reg_space[5620] = 8'h00;
reg_space[5621] = 8'h00;
reg_space[5622] = 8'h00;
reg_space[5623] = 8'h00;
reg_space[5624] = 8'h00;
reg_space[5625] = 8'h00;
reg_space[5626] = 8'h00;
reg_space[5627] = 8'h00;
reg_space[5628] = 8'h00;
reg_space[5629] = 8'h00;
reg_space[5630] = 8'h00;
reg_space[5631] = 8'h00;
reg_space[5632] = 8'h00;
reg_space[5633] = 8'h00;
reg_space[5634] = 8'h00;
reg_space[5635] = 8'h00;
reg_space[5636] = 8'h00;
reg_space[5637] = 8'h00;
reg_space[5638] = 8'h00;
reg_space[5639] = 8'h00;
reg_space[5640] = 8'h00;
reg_space[5641] = 8'h00;
reg_space[5642] = 8'h00;
reg_space[5643] = 8'h00;
reg_space[5644] = 8'h00;
reg_space[5645] = 8'h00;
reg_space[5646] = 8'h00;
reg_space[5647] = 8'h00;
reg_space[5648] = 8'h00;
reg_space[5649] = 8'h00;
reg_space[5650] = 8'h00;
reg_space[5651] = 8'h00;
reg_space[5652] = 8'h00;
reg_space[5653] = 8'h00;
reg_space[5654] = 8'h00;
reg_space[5655] = 8'h00;
reg_space[5656] = 8'h00;
reg_space[5657] = 8'h00;
reg_space[5658] = 8'h00;
reg_space[5659] = 8'h00;
reg_space[5660] = 8'h00;
reg_space[5661] = 8'h00;
reg_space[5662] = 8'h00;
reg_space[5663] = 8'h00;
reg_space[5664] = 8'h00;
reg_space[5665] = 8'h00;
reg_space[5666] = 8'h00;
reg_space[5667] = 8'h00;
reg_space[5668] = 8'h00;
reg_space[5669] = 8'h00;
reg_space[5670] = 8'h00;
reg_space[5671] = 8'h00;
reg_space[5672] = 8'h00;
reg_space[5673] = 8'h00;
reg_space[5674] = 8'h00;
reg_space[5675] = 8'h00;
reg_space[5676] = 8'h00;
reg_space[5677] = 8'h00;
reg_space[5678] = 8'h00;
reg_space[5679] = 8'h00;
reg_space[5680] = 8'h00;
reg_space[5681] = 8'h00;
reg_space[5682] = 8'h00;
reg_space[5683] = 8'h00;
reg_space[5684] = 8'h00;
reg_space[5685] = 8'h00;
reg_space[5686] = 8'h00;
reg_space[5687] = 8'h00;
reg_space[5688] = 8'h00;
reg_space[5689] = 8'h00;
reg_space[5690] = 8'h00;
reg_space[5691] = 8'h00;
reg_space[5692] = 8'h00;
reg_space[5693] = 8'h00;
reg_space[5694] = 8'h00;
reg_space[5695] = 8'h00;
reg_space[5696] = 8'h00;
reg_space[5697] = 8'h00;
reg_space[5698] = 8'h00;
reg_space[5699] = 8'h00;
reg_space[5700; = 8'h00;
reg_space[5701] = 8'h00;
reg_space[5702] = 8'h00;
reg_space[5703] = 8'h00;
reg_space[5704] = 8'h00;
reg_space[5705] = 8'h00;
reg_space[5706] = 8'h00;
reg_space[5707] = 8'h00;
reg_space[5708] = 8'h00;
reg_space[5709] = 8'h00;
reg_space[5710] = 8'h00;
reg_space[5711] = 8'h00;
reg_space[5712] = 8'h00;
reg_space[5713] = 8'h00;
reg_space[5714] = 8'h00;
reg_space[5715] = 8'h00;
reg_space[5716] = 8'h00;
reg_space[5717] = 8'h00;
reg_space[5718] = 8'h00;
reg_space[5719] = 8'h00;
reg_space[5720] = 8'h00;
reg_space[5721] = 8'h00;
reg_space[5722] = 8'h00;
reg_space[5723] = 8'h00;
reg_space[5724] = 8'h00;
reg_space[5725] = 8'h00;
reg_space[5726] = 8'h00;
reg_space[5727] = 8'h00;
reg_space[5728] = 8'h00;
reg_space[5729] = 8'h00;
reg_space[5730] = 8'h00;
reg_space[5731] = 8'h00;
reg_space[5732] = 8'h00;
reg_space[5733] = 8'h00;
reg_space[5734] = 8'h00;
reg_space[5735] = 8'h00;
reg_space[5736] = 8'h00;
reg_space[5737] = 8'h00;
reg_space[5738] = 8'h00;
reg_space[5739] = 8'h00;
reg_space[5740] = 8'h00;
reg_space[5741] = 8'h00;
reg_space[5742] = 8'h00;
reg_space[5743] = 8'h00;
reg_space[5744] = 8'h00;
reg_space[5745] = 8'h00;
reg_space[5746] = 8'h00;
reg_space[5747] = 8'h00;
reg_space[5748] = 8'h00;
reg_space[5749] = 8'h00;
reg_space[5750] = 8'h00;
reg_space[5751] = 8'h00;
reg_space[5752] = 8'h00;
reg_space[5753] = 8'h00;
reg_space[5754] = 8'h00;
reg_space[5755] = 8'h00;
reg_space[5756] = 8'h00;
reg_space[5757] = 8'h00;
reg_space[5758] = 8'h00;
reg_space[5759] = 8'h00;
reg_space[5760] = 8'h00;
reg_space[5761] = 8'h00;
reg_space[5762] = 8'h00;
reg_space[5763] = 8'h00;
reg_space[5764] = 8'h00;
reg_space[5765] = 8'h00;
reg_space[5766] = 8'h00;
reg_space[5767] = 8'h00;
reg_space[5768] = 8'h00;
reg_space[5769] = 8'h00;
reg_space[5770] = 8'h00;
reg_space[5771] = 8'h00;
reg_space[5772] = 8'h00;
reg_space[5773] = 8'h00;
reg_space[5774] = 8'h00;
reg_space[5775] = 8'h00;
reg_space[5776] = 8'h00;
reg_space[5777] = 8'h00;
reg_space[5778] = 8'h00;
reg_space[5779] = 8'h00;
reg_space[5780] = 8'h00;
reg_space[5781] = 8'h00;
reg_space[5782] = 8'h00;
reg_space[5783] = 8'h00;
reg_space[5784] = 8'h00;
reg_space[5785] = 8'h00;
reg_space[5786] = 8'h00;
reg_space[5787] = 8'h00;
reg_space[5788] = 8'h00;
reg_space[5789] = 8'h00;
reg_space[5790] = 8'h00;
reg_space[5791] = 8'h00;
reg_space[5792] = 8'h00;
reg_space[5793] = 8'h00;
reg_space[5794] = 8'h00;
reg_space[5795] = 8'h00;
reg_space[5796] = 8'h00;
reg_space[5797] = 8'h00;
reg_space[5798] = 8'h00;
reg_space[5799] = 8'h00;
reg_space[5800; = 8'h00;
reg_space[5801] = 8'h00;
reg_space[5802] = 8'h00;
reg_space[5803] = 8'h00;
reg_space[5804] = 8'h00;
reg_space[5805] = 8'h00;
reg_space[5806] = 8'h00;
reg_space[5807] = 8'h00;
reg_space[5808] = 8'h00;
reg_space[5809] = 8'h00;
reg_space[5810] = 8'h00;
reg_space[5811] = 8'h00;
reg_space[5812] = 8'h00;
reg_space[5813] = 8'h00;
reg_space[5814] = 8'h00;
reg_space[5815] = 8'h00;
reg_space[5816] = 8'h00;
reg_space[5817] = 8'h00;
reg_space[5818] = 8'h00;
reg_space[5819] = 8'h00;
reg_space[5820] = 8'h00;
reg_space[5821] = 8'h00;
reg_space[5822] = 8'h00;
reg_space[5823] = 8'h00;
reg_space[5824] = 8'h00;
reg_space[5825] = 8'h00;
reg_space[5826] = 8'h00;
reg_space[5827] = 8'h00;
reg_space[5828] = 8'h00;
reg_space[5829] = 8'h00;
reg_space[5830] = 8'h00;
reg_space[5831] = 8'h00;
reg_space[5832] = 8'h00;
reg_space[5833] = 8'h00;
reg_space[5834] = 8'h00;
reg_space[5835] = 8'h00;
reg_space[5836] = 8'h00;
reg_space[5837] = 8'h00;
reg_space[5838] = 8'h00;
reg_space[5839] = 8'h00;
reg_space[5840] = 8'h00;
reg_space[5841] = 8'h00;
reg_space[5842] = 8'h00;
reg_space[5843] = 8'h00;
reg_space[5844] = 8'h00;
reg_space[5845] = 8'h00;
reg_space[5846] = 8'h00;
reg_space[5847] = 8'h00;
reg_space[5848] = 8'h00;
reg_space[5849] = 8'h00;
reg_space[5850] = 8'h00;
reg_space[5851] = 8'h00;
reg_space[5852] = 8'h00;
reg_space[5853] = 8'h00;
reg_space[5854] = 8'h00;
reg_space[5855] = 8'h00;
reg_space[5856] = 8'h00;
reg_space[5857] = 8'h00;
reg_space[5858] = 8'h00;
reg_space[5859] = 8'h00;
reg_space[5860] = 8'h00;
reg_space[5861] = 8'h00;
reg_space[5862] = 8'h00;
reg_space[5863] = 8'h00;
reg_space[5864] = 8'h00;
reg_space[5865] = 8'h00;
reg_space[5866] = 8'h00;
reg_space[5867] = 8'h00;
reg_space[5868] = 8'h00;
reg_space[5869] = 8'h00;
reg_space[5870] = 8'h00;
reg_space[5871] = 8'h00;
reg_space[5872] = 8'h00;
reg_space[5873] = 8'h00;
reg_space[5874] = 8'h00;
reg_space[5875] = 8'h00;
reg_space[5876] = 8'h00;
reg_space[5877] = 8'h00;
reg_space[5878] = 8'h00;
reg_space[5879] = 8'h00;
reg_space[5880] = 8'h00;
reg_space[5881] = 8'h00;
reg_space[5882] = 8'h00;
reg_space[5883] = 8'h00;
reg_space[5884] = 8'h00;
reg_space[5885] = 8'h00;
reg_space[5886] = 8'h00;
reg_space[5887] = 8'h00;
reg_space[5888] = 8'h00;
reg_space[5889] = 8'h00;
reg_space[5890] = 8'h00;
reg_space[5891] = 8'h00;
reg_space[5892] = 8'h00;
reg_space[5893] = 8'h00;
reg_space[5894] = 8'h00;
reg_space[5895] = 8'h00;
reg_space[5896] = 8'h00;
reg_space[5897] = 8'h00;
reg_space[5898] = 8'h00;
reg_space[5899] = 8'h00;
reg_space[5900; = 8'h00;
reg_space[5901] = 8'h00;
reg_space[5902] = 8'h00;
reg_space[5903] = 8'h00;
reg_space[5904] = 8'h00;
reg_space[5905] = 8'h00;
reg_space[5906] = 8'h00;
reg_space[5907] = 8'h00;
reg_space[5908] = 8'h00;
reg_space[5909] = 8'h00;
reg_space[5910] = 8'h00;
reg_space[5911] = 8'h00;
reg_space[5912] = 8'h00;
reg_space[5913] = 8'h00;
reg_space[5914] = 8'h00;
reg_space[5915] = 8'h00;
reg_space[5916] = 8'h00;
reg_space[5917] = 8'h00;
reg_space[5918] = 8'h00;
reg_space[5919] = 8'h00;
reg_space[5920] = 8'h00;
reg_space[5921] = 8'h00;
reg_space[5922] = 8'h00;
reg_space[5923] = 8'h00;
reg_space[5924] = 8'h00;
reg_space[5925] = 8'h00;
reg_space[5926] = 8'h00;
reg_space[5927] = 8'h00;
reg_space[5928] = 8'h00;
reg_space[5929] = 8'h00;
reg_space[5930] = 8'h00;
reg_space[5931] = 8'h00;
reg_space[5932] = 8'h00;
reg_space[5933] = 8'h00;
reg_space[5934] = 8'h00;
reg_space[5935] = 8'h00;
reg_space[5936] = 8'h00;
reg_space[5937] = 8'h00;
reg_space[5938] = 8'h00;
reg_space[5939] = 8'h00;
reg_space[5940] = 8'h00;
reg_space[5941] = 8'h00;
reg_space[5942] = 8'h00;
reg_space[5943] = 8'h00;
reg_space[5944] = 8'h00;
reg_space[5945] = 8'h00;
reg_space[5946] = 8'h00;
reg_space[5947] = 8'h00;
reg_space[5948] = 8'h00;
reg_space[5949] = 8'h00;
reg_space[5950] = 8'h00;
reg_space[5951] = 8'h00;
reg_space[5952] = 8'h00;
reg_space[5953] = 8'h00;
reg_space[5954] = 8'h00;
reg_space[5955] = 8'h00;
reg_space[5956] = 8'h00;
reg_space[5957] = 8'h00;
reg_space[5958] = 8'h00;
reg_space[5959] = 8'h00;
reg_space[5960] = 8'h00;
reg_space[5961] = 8'h00;
reg_space[5962] = 8'h00;
reg_space[5963] = 8'h00;
reg_space[5964] = 8'h00;
reg_space[5965] = 8'h00;
reg_space[5966] = 8'h00;
reg_space[5967] = 8'h00;
reg_space[5968] = 8'h00;
reg_space[5969] = 8'h00;
reg_space[5970] = 8'h00;
reg_space[5971] = 8'h00;
reg_space[5972] = 8'h00;
reg_space[5973] = 8'h00;
reg_space[5974] = 8'h00;
reg_space[5975] = 8'h00;
reg_space[5976] = 8'h00;
reg_space[5977] = 8'h00;
reg_space[5978] = 8'h00;
reg_space[5979] = 8'h00;
reg_space[5980] = 8'h00;
reg_space[5981] = 8'h00;
reg_space[5982] = 8'h00;
reg_space[5983] = 8'h00;
reg_space[5984] = 8'h00;
reg_space[5985] = 8'h00;
reg_space[5986] = 8'h00;
reg_space[5987] = 8'h00;
reg_space[5988] = 8'h00;
reg_space[5989] = 8'h00;
reg_space[5990] = 8'h00;
reg_space[5991] = 8'h00;
reg_space[5992] = 8'h00;
reg_space[5993] = 8'h00;
reg_space[5994] = 8'h00;
reg_space[5995] = 8'h00;
reg_space[5996] = 8'h00;
reg_space[5997] = 8'h00;
reg_space[5998] = 8'h00;
reg_space[5999] = 8'h00;
reg_space[600;0] = 8'h00;
reg_space[600;1] = 8'h00;
reg_space[600;2] = 8'h00;
reg_space[600;3] = 8'h00;
reg_space[600;4] = 8'h00;
reg_space[600;5] = 8'h00;
reg_space[600;6] = 8'h00;
reg_space[600;7] = 8'h00;
reg_space[600;8] = 8'h00;
reg_space[600;9] = 8'h00;
reg_space[6010] = 8'h00;
reg_space[6011] = 8'h00;
reg_space[6012] = 8'h00;
reg_space[6013] = 8'h00;
reg_space[6014] = 8'h00;
reg_space[6015] = 8'h00;
reg_space[6016] = 8'h00;
reg_space[6017] = 8'h00;
reg_space[6018] = 8'h00;
reg_space[6019] = 8'h00;
reg_space[6020] = 8'h00;
reg_space[6021] = 8'h00;
reg_space[6022] = 8'h00;
reg_space[6023] = 8'h00;
reg_space[6024] = 8'h00;
reg_space[6025] = 8'h00;
reg_space[6026] = 8'h00;
reg_space[6027] = 8'h00;
reg_space[6028] = 8'h00;
reg_space[6029] = 8'h00;
reg_space[6030] = 8'h00;
reg_space[6031] = 8'h00;
reg_space[6032] = 8'h00;
reg_space[6033] = 8'h00;
reg_space[6034] = 8'h00;
reg_space[6035] = 8'h00;
reg_space[6036] = 8'h00;
reg_space[6037] = 8'h00;
reg_space[6038] = 8'h00;
reg_space[6039] = 8'h00;
reg_space[6040] = 8'h00;
reg_space[6041] = 8'h00;
reg_space[6042] = 8'h00;
reg_space[6043] = 8'h00;
reg_space[6044] = 8'h00;
reg_space[6045] = 8'h00;
reg_space[6046] = 8'h00;
reg_space[6047] = 8'h00;
reg_space[6048] = 8'h00;
reg_space[6049] = 8'h00;
reg_space[6050] = 8'h00;
reg_space[6051] = 8'h00;
reg_space[6052] = 8'h00;
reg_space[6053] = 8'h00;
reg_space[6054] = 8'h00;
reg_space[6055] = 8'h00;
reg_space[6056] = 8'h00;
reg_space[6057] = 8'h00;
reg_space[6058] = 8'h00;
reg_space[6059] = 8'h00;
reg_space[6060] = 8'h00;
reg_space[6061] = 8'h00;
reg_space[6062] = 8'h00;
reg_space[6063] = 8'h00;
reg_space[6064] = 8'h00;
reg_space[6065] = 8'h00;
reg_space[6066] = 8'h00;
reg_space[6067] = 8'h00;
reg_space[6068] = 8'h00;
reg_space[6069] = 8'h00;
reg_space[6070] = 8'h00;
reg_space[6071] = 8'h00;
reg_space[6072] = 8'h00;
reg_space[6073] = 8'h00;
reg_space[6074] = 8'h00;
reg_space[6075] = 8'h00;
reg_space[6076] = 8'h00;
reg_space[6077] = 8'h00;
reg_space[6078] = 8'h00;
reg_space[6079] = 8'h00;
reg_space[6080] = 8'h00;
reg_space[6081] = 8'h00;
reg_space[6082] = 8'h00;
reg_space[6083] = 8'h00;
reg_space[6084] = 8'h00;
reg_space[6085] = 8'h00;
reg_space[6086] = 8'h00;
reg_space[6087] = 8'h00;
reg_space[6088] = 8'h00;
reg_space[6089] = 8'h00;
reg_space[6090] = 8'h00;
reg_space[6091] = 8'h00;
reg_space[6092] = 8'h00;
reg_space[6093] = 8'h00;
reg_space[6094] = 8'h00;
reg_space[6095] = 8'h00;
reg_space[6096] = 8'h00;
reg_space[6097] = 8'h00;
reg_space[6098] = 8'h00;
reg_space[6099] = 8'h00;
reg_space[6100; = 8'h00;
reg_space[6101] = 8'h00;
reg_space[6102] = 8'h00;
reg_space[6103] = 8'h00;
reg_space[6104] = 8'h00;
reg_space[6105] = 8'h00;
reg_space[6106] = 8'h00;
reg_space[6107] = 8'h00;
reg_space[6108] = 8'h00;
reg_space[6109] = 8'h00;
reg_space[6110] = 8'h00;
reg_space[6111] = 8'h00;
reg_space[6112] = 8'h00;
reg_space[6113] = 8'h00;
reg_space[6114] = 8'h00;
reg_space[6115] = 8'h00;
reg_space[6116] = 8'h00;
reg_space[6117] = 8'h00;
reg_space[6118] = 8'h00;
reg_space[6119] = 8'h00;
reg_space[6120] = 8'h00;
reg_space[6121] = 8'h00;
reg_space[6122] = 8'h00;
reg_space[6123] = 8'h00;
reg_space[6124] = 8'h00;
reg_space[6125] = 8'h00;
reg_space[6126] = 8'h00;
reg_space[6127] = 8'h00;
reg_space[6128] = 8'h00;
reg_space[6129] = 8'h00;
reg_space[6130] = 8'h00;
reg_space[6131] = 8'h00;
reg_space[6132] = 8'h00;
reg_space[6133] = 8'h00;
reg_space[6134] = 8'h00;
reg_space[6135] = 8'h00;
reg_space[6136] = 8'h00;
reg_space[6137] = 8'h00;
reg_space[6138] = 8'h00;
reg_space[6139] = 8'h00;
reg_space[6140] = 8'h00;
reg_space[6141] = 8'h00;
reg_space[6142] = 8'h00;
reg_space[6143] = 8'h00;
reg_space[6144] = 8'h00;
reg_space[6145] = 8'h00;
reg_space[6146] = 8'h00;
reg_space[6147] = 8'h00;
reg_space[6148] = 8'h00;
reg_space[6149] = 8'h00;
reg_space[6150] = 8'h00;
reg_space[6151] = 8'h00;
reg_space[6152] = 8'h00;
reg_space[6153] = 8'h00;
reg_space[6154] = 8'h00;
reg_space[6155] = 8'h00;
reg_space[6156] = 8'h00;
reg_space[6157] = 8'h00;
reg_space[6158] = 8'h00;
reg_space[6159] = 8'h00;
reg_space[6160] = 8'h00;
reg_space[6161] = 8'h00;
reg_space[6162] = 8'h00;
reg_space[6163] = 8'h00;
reg_space[6164] = 8'h00;
reg_space[6165] = 8'h00;
reg_space[6166] = 8'h00;
reg_space[6167] = 8'h00;
reg_space[6168] = 8'h00;
reg_space[6169] = 8'h00;
reg_space[6170] = 8'h00;
reg_space[6171] = 8'h00;
reg_space[6172] = 8'h00;
reg_space[6173] = 8'h00;
reg_space[6174] = 8'h00;
reg_space[6175] = 8'h00;
reg_space[6176] = 8'h00;
reg_space[6177] = 8'h00;
reg_space[6178] = 8'h00;
reg_space[6179] = 8'h00;
reg_space[6180] = 8'h00;
reg_space[6181] = 8'h00;
reg_space[6182] = 8'h00;
reg_space[6183] = 8'h00;
reg_space[6184] = 8'h00;
reg_space[6185] = 8'h00;
reg_space[6186] = 8'h00;
reg_space[6187] = 8'h00;
reg_space[6188] = 8'h00;
reg_space[6189] = 8'h00;
reg_space[6190] = 8'h00;
reg_space[6191] = 8'h00;
reg_space[6192] = 8'h00;
reg_space[6193] = 8'h00;
reg_space[6194] = 8'h00;
reg_space[6195] = 8'h00;
reg_space[6196] = 8'h00;
reg_space[6197] = 8'h00;
reg_space[6198] = 8'h00;
reg_space[6199] = 8'h00;
reg_space[6200; = 8'h00;
reg_space[6201] = 8'h00;
reg_space[6202] = 8'h00;
reg_space[6203] = 8'h00;
reg_space[6204] = 8'h00;
reg_space[6205] = 8'h00;
reg_space[6206] = 8'h00;
reg_space[6207] = 8'h00;
reg_space[6208] = 8'h00;
reg_space[6209] = 8'h00;
reg_space[6210] = 8'h00;
reg_space[6211] = 8'h00;
reg_space[6212] = 8'h00;
reg_space[6213] = 8'h00;
reg_space[6214] = 8'h00;
reg_space[6215] = 8'h00;
reg_space[6216] = 8'h00;
reg_space[6217] = 8'h00;
reg_space[6218] = 8'h00;
reg_space[6219] = 8'h00;
reg_space[6220] = 8'h00;
reg_space[6221] = 8'h00;
reg_space[6222] = 8'h00;
reg_space[6223] = 8'h00;
reg_space[6224] = 8'h00;
reg_space[6225] = 8'h00;
reg_space[6226] = 8'h00;
reg_space[6227] = 8'h00;
reg_space[6228] = 8'h00;
reg_space[6229] = 8'h00;
reg_space[6230] = 8'h00;
reg_space[6231] = 8'h00;
reg_space[6232] = 8'h00;
reg_space[6233] = 8'h00;
reg_space[6234] = 8'h00;
reg_space[6235] = 8'h00;
reg_space[6236] = 8'h00;
reg_space[6237] = 8'h00;
reg_space[6238] = 8'h00;
reg_space[6239] = 8'h00;
reg_space[6240] = 8'h00;
reg_space[6241] = 8'h00;
reg_space[6242] = 8'h00;
reg_space[6243] = 8'h00;
reg_space[6244] = 8'h00;
reg_space[6245] = 8'h00;
reg_space[6246] = 8'h00;
reg_space[6247] = 8'h00;
reg_space[6248] = 8'h00;
reg_space[6249] = 8'h00;
reg_space[6250] = 8'h00;
reg_space[6251] = 8'h00;
reg_space[6252] = 8'h00;
reg_space[6253] = 8'h00;
reg_space[6254] = 8'h00;
reg_space[6255] = 8'h00;
reg_space[6256] = 8'h00;
reg_space[6257] = 8'h00;
reg_space[6258] = 8'h00;
reg_space[6259] = 8'h00;
reg_space[6260] = 8'h00;
reg_space[6261] = 8'h00;
reg_space[6262] = 8'h00;
reg_space[6263] = 8'h00;
reg_space[6264] = 8'h00;
reg_space[6265] = 8'h00;
reg_space[6266] = 8'h00;
reg_space[6267] = 8'h00;
reg_space[6268] = 8'h00;
reg_space[6269] = 8'h00;
reg_space[6270] = 8'h00;
reg_space[6271] = 8'h00;
reg_space[6272] = 8'h00;
reg_space[6273] = 8'h00;
reg_space[6274] = 8'h00;
reg_space[6275] = 8'h00;
reg_space[6276] = 8'h00;
reg_space[6277] = 8'h00;
reg_space[6278] = 8'h00;
reg_space[6279] = 8'h00;
reg_space[6280] = 8'h00;
reg_space[6281] = 8'h00;
reg_space[6282] = 8'h00;
reg_space[6283] = 8'h00;
reg_space[6284] = 8'h00;
reg_space[6285] = 8'h00;
reg_space[6286] = 8'h00;
reg_space[6287] = 8'h00;
reg_space[6288] = 8'h00;
reg_space[6289] = 8'h00;
reg_space[6290] = 8'h00;
reg_space[6291] = 8'h00;
reg_space[6292] = 8'h00;
reg_space[6293] = 8'h00;
reg_space[6294] = 8'h00;
reg_space[6295] = 8'h00;
reg_space[6296] = 8'h00;
reg_space[6297] = 8'h00;
reg_space[6298] = 8'h00;
reg_space[6299] = 8'h00;
reg_space[6300; = 8'h00;
reg_space[6301] = 8'h00;
reg_space[6302] = 8'h00;
reg_space[6303] = 8'h00;
reg_space[6304] = 8'h00;
reg_space[6305] = 8'h00;
reg_space[6306] = 8'h00;
reg_space[6307] = 8'h00;
reg_space[6308] = 8'h00;
reg_space[6309] = 8'h00;
reg_space[6310] = 8'h00;
reg_space[6311] = 8'h00;
reg_space[6312] = 8'h00;
reg_space[6313] = 8'h00;
reg_space[6314] = 8'h00;
reg_space[6315] = 8'h00;
reg_space[6316] = 8'h00;
reg_space[6317] = 8'h00;
reg_space[6318] = 8'h00;
reg_space[6319] = 8'h00;
reg_space[6320] = 8'h00;
reg_space[6321] = 8'h00;
reg_space[6322] = 8'h00;
reg_space[6323] = 8'h00;
reg_space[6324] = 8'h00;
reg_space[6325] = 8'h00;
reg_space[6326] = 8'h00;
reg_space[6327] = 8'h00;
reg_space[6328] = 8'h00;
reg_space[6329] = 8'h00;
reg_space[6330] = 8'h00;
reg_space[6331] = 8'h00;
reg_space[6332] = 8'h00;
reg_space[6333] = 8'h00;
reg_space[6334] = 8'h00;
reg_space[6335] = 8'h00;
reg_space[6336] = 8'h00;
reg_space[6337] = 8'h00;
reg_space[6338] = 8'h00;
reg_space[6339] = 8'h00;
reg_space[6340] = 8'h00;
reg_space[6341] = 8'h00;
reg_space[6342] = 8'h00;
reg_space[6343] = 8'h00;
reg_space[6344] = 8'h00;
reg_space[6345] = 8'h00;
reg_space[6346] = 8'h00;
reg_space[6347] = 8'h00;
reg_space[6348] = 8'h00;
reg_space[6349] = 8'h00;
reg_space[6350] = 8'h00;
reg_space[6351] = 8'h00;
reg_space[6352] = 8'h00;
reg_space[6353] = 8'h00;
reg_space[6354] = 8'h00;
reg_space[6355] = 8'h00;
reg_space[6356] = 8'h00;
reg_space[6357] = 8'h00;
reg_space[6358] = 8'h00;
reg_space[6359] = 8'h00;
reg_space[6360] = 8'h00;
reg_space[6361] = 8'h00;
reg_space[6362] = 8'h00;
reg_space[6363] = 8'h00;
reg_space[6364] = 8'h00;
reg_space[6365] = 8'h00;
reg_space[6366] = 8'h00;
reg_space[6367] = 8'h00;
reg_space[6368] = 8'h00;
reg_space[6369] = 8'h00;
reg_space[6370] = 8'h00;
reg_space[6371] = 8'h00;
reg_space[6372] = 8'h00;
reg_space[6373] = 8'h00;
reg_space[6374] = 8'h00;
reg_space[6375] = 8'h00;
reg_space[6376] = 8'h00;
reg_space[6377] = 8'h00;
reg_space[6378] = 8'h00;
reg_space[6379] = 8'h00;
reg_space[6380] = 8'h00;
reg_space[6381] = 8'h00;
reg_space[6382] = 8'h00;
reg_space[6383] = 8'h00;
reg_space[6384] = 8'h00;
reg_space[6385] = 8'h00;
reg_space[6386] = 8'h00;
reg_space[6387] = 8'h00;
reg_space[6388] = 8'h00;
reg_space[6389] = 8'h00;
reg_space[6390] = 8'h00;
reg_space[6391] = 8'h00;
reg_space[6392] = 8'h00;
reg_space[6393] = 8'h00;
reg_space[6394] = 8'h00;
reg_space[6395] = 8'h00;
reg_space[6396] = 8'h00;
reg_space[6397] = 8'h00;
reg_space[6398] = 8'h00;
reg_space[6399] = 8'h00;
reg_space[6400; = 8'h00;
reg_space[6401] = 8'h00;
reg_space[6402] = 8'h00;
reg_space[6403] = 8'h00;
reg_space[6404] = 8'h00;
reg_space[6405] = 8'h00;
reg_space[6406] = 8'h00;
reg_space[6407] = 8'h00;
reg_space[6408] = 8'h00;
reg_space[6409] = 8'h00;
reg_space[6410] = 8'h00;
reg_space[6411] = 8'h00;
reg_space[6412] = 8'h00;
reg_space[6413] = 8'h00;
reg_space[6414] = 8'h00;
reg_space[6415] = 8'h00;
reg_space[6416] = 8'h00;
reg_space[6417] = 8'h00;
reg_space[6418] = 8'h00;
reg_space[6419] = 8'h00;
reg_space[6420] = 8'h00;
reg_space[6421] = 8'h00;
reg_space[6422] = 8'h00;
reg_space[6423] = 8'h00;
reg_space[6424] = 8'h00;
reg_space[6425] = 8'h00;
reg_space[6426] = 8'h00;
reg_space[6427] = 8'h00;
reg_space[6428] = 8'h00;
reg_space[6429] = 8'h00;
reg_space[6430] = 8'h00;
reg_space[6431] = 8'h00;
reg_space[6432] = 8'h00;
reg_space[6433] = 8'h00;
reg_space[6434] = 8'h00;
reg_space[6435] = 8'h00;
reg_space[6436] = 8'h00;
reg_space[6437] = 8'h00;
reg_space[6438] = 8'h00;
reg_space[6439] = 8'h00;
reg_space[6440] = 8'h00;
reg_space[6441] = 8'h00;
reg_space[6442] = 8'h00;
reg_space[6443] = 8'h00;
reg_space[6444] = 8'h00;
reg_space[6445] = 8'h00;
reg_space[6446] = 8'h00;
reg_space[6447] = 8'h00;
reg_space[6448] = 8'h00;
reg_space[6449] = 8'h00;
reg_space[6450] = 8'h00;
reg_space[6451] = 8'h00;
reg_space[6452] = 8'h00;
reg_space[6453] = 8'h00;
reg_space[6454] = 8'h00;
reg_space[6455] = 8'h00;
reg_space[6456] = 8'h00;
reg_space[6457] = 8'h00;
reg_space[6458] = 8'h00;
reg_space[6459] = 8'h00;
reg_space[6460] = 8'h00;
reg_space[6461] = 8'h00;
reg_space[6462] = 8'h00;
reg_space[6463] = 8'h00;
reg_space[6464] = 8'h00;
reg_space[6465] = 8'h00;
reg_space[6466] = 8'h00;
reg_space[6467] = 8'h00;
reg_space[6468] = 8'h00;
reg_space[6469] = 8'h00;
reg_space[6470] = 8'h00;
reg_space[6471] = 8'h00;
reg_space[6472] = 8'h00;
reg_space[6473] = 8'h00;
reg_space[6474] = 8'h00;
reg_space[6475] = 8'h00;
reg_space[6476] = 8'h00;
reg_space[6477] = 8'h00;
reg_space[6478] = 8'h00;
reg_space[6479] = 8'h00;
reg_space[6480] = 8'h00;
reg_space[6481] = 8'h00;
reg_space[6482] = 8'h00;
reg_space[6483] = 8'h00;
reg_space[6484] = 8'h00;
reg_space[6485] = 8'h00;
reg_space[6486] = 8'h00;
reg_space[6487] = 8'h00;
reg_space[6488] = 8'h00;
reg_space[6489] = 8'h00;
reg_space[6490] = 8'h00;
reg_space[6491] = 8'h00;
reg_space[6492] = 8'h00;
reg_space[6493] = 8'h00;
reg_space[6494] = 8'h00;
reg_space[6495] = 8'h00;
reg_space[6496] = 8'h00;
reg_space[6497] = 8'h00;
reg_space[6498] = 8'h00;
reg_space[6499] = 8'h00;
reg_space[6500; = 8'h00;
reg_space[6501] = 8'h00;
reg_space[6502] = 8'h00;
reg_space[6503] = 8'h00;
reg_space[6504] = 8'h00;
reg_space[6505] = 8'h00;
reg_space[6506] = 8'h00;
reg_space[6507] = 8'h00;
reg_space[6508] = 8'h00;
reg_space[6509] = 8'h00;
reg_space[6510] = 8'h00;
reg_space[6511] = 8'h00;
reg_space[6512] = 8'h00;
reg_space[6513] = 8'h00;
reg_space[6514] = 8'h00;
reg_space[6515] = 8'h00;
reg_space[6516] = 8'h00;
reg_space[6517] = 8'h00;
reg_space[6518] = 8'h00;
reg_space[6519] = 8'h00;
reg_space[6520] = 8'h00;
reg_space[6521] = 8'h00;
reg_space[6522] = 8'h00;
reg_space[6523] = 8'h00;
reg_space[6524] = 8'h00;
reg_space[6525] = 8'h00;
reg_space[6526] = 8'h00;
reg_space[6527] = 8'h00;
reg_space[6528] = 8'h00;
reg_space[6529] = 8'h00;
reg_space[6530] = 8'h00;
reg_space[6531] = 8'h00;
reg_space[6532] = 8'h00;
reg_space[6533] = 8'h00;
reg_space[6534] = 8'h00;
reg_space[6535] = 8'h00;
reg_space[6536] = 8'h00;
reg_space[6537] = 8'h00;
reg_space[6538] = 8'h00;
reg_space[6539] = 8'h00;
reg_space[6540] = 8'h00;
reg_space[6541] = 8'h00;
reg_space[6542] = 8'h00;
reg_space[6543] = 8'h00;
reg_space[6544] = 8'h00;
reg_space[6545] = 8'h00;
reg_space[6546] = 8'h00;
reg_space[6547] = 8'h00;
reg_space[6548] = 8'h00;
reg_space[6549] = 8'h00;
reg_space[6550] = 8'h00;
reg_space[6551] = 8'h00;
reg_space[6552] = 8'h00;
reg_space[6553] = 8'h00;
reg_space[6554] = 8'h00;
reg_space[6555] = 8'h00;
reg_space[6556] = 8'h00;
reg_space[6557] = 8'h00;
reg_space[6558] = 8'h00;
reg_space[6559] = 8'h00;
reg_space[6560] = 8'h00;
reg_space[6561] = 8'h00;
reg_space[6562] = 8'h00;
reg_space[6563] = 8'h00;
reg_space[6564] = 8'h00;
reg_space[6565] = 8'h00;
reg_space[6566] = 8'h00;
reg_space[6567] = 8'h00;
reg_space[6568] = 8'h00;
reg_space[6569] = 8'h00;
reg_space[6570] = 8'h00;
reg_space[6571] = 8'h00;
reg_space[6572] = 8'h00;
reg_space[6573] = 8'h00;
reg_space[6574] = 8'h00;
reg_space[6575] = 8'h00;
reg_space[6576] = 8'h00;
reg_space[6577] = 8'h00;
reg_space[6578] = 8'h00;
reg_space[6579] = 8'h00;
reg_space[6580] = 8'h00;
reg_space[6581] = 8'h00;
reg_space[6582] = 8'h00;
reg_space[6583] = 8'h00;
reg_space[6584] = 8'h00;
reg_space[6585] = 8'h00;
reg_space[6586] = 8'h00;
reg_space[6587] = 8'h00;
reg_space[6588] = 8'h00;
reg_space[6589] = 8'h00;
reg_space[6590] = 8'h00;
reg_space[6591] = 8'h00;
reg_space[6592] = 8'h00;
reg_space[6593] = 8'h00;
reg_space[6594] = 8'h00;
reg_space[6595] = 8'h00;
reg_space[6596] = 8'h00;
reg_space[6597] = 8'h00;
reg_space[6598] = 8'h00;
reg_space[6599] = 8'h00;
reg_space[6600; = 8'h00;
reg_space[6601] = 8'h00;
reg_space[6602] = 8'h00;
reg_space[6603] = 8'h00;
reg_space[6604] = 8'h00;
reg_space[6605] = 8'h00;
reg_space[6606] = 8'h00;
reg_space[6607] = 8'h00;
reg_space[6608] = 8'h00;
reg_space[6609] = 8'h00;
reg_space[6610] = 8'h00;
reg_space[6611] = 8'h00;
reg_space[6612] = 8'h00;
reg_space[6613] = 8'h00;
reg_space[6614] = 8'h00;
reg_space[6615] = 8'h00;
reg_space[6616] = 8'h00;
reg_space[6617] = 8'h00;
reg_space[6618] = 8'h00;
reg_space[6619] = 8'h00;
reg_space[6620] = 8'h00;
reg_space[6621] = 8'h00;
reg_space[6622] = 8'h00;
reg_space[6623] = 8'h00;
reg_space[6624] = 8'h00;
reg_space[6625] = 8'h00;
reg_space[6626] = 8'h00;
reg_space[6627] = 8'h00;
reg_space[6628] = 8'h00;
reg_space[6629] = 8'h00;
reg_space[6630] = 8'h00;
reg_space[6631] = 8'h00;
reg_space[6632] = 8'h00;
reg_space[6633] = 8'h00;
reg_space[6634] = 8'h00;
reg_space[6635] = 8'h00;
reg_space[6636] = 8'h00;
reg_space[6637] = 8'h00;
reg_space[6638] = 8'h00;
reg_space[6639] = 8'h00;
reg_space[6640] = 8'h00;
reg_space[6641] = 8'h00;
reg_space[6642] = 8'h00;
reg_space[6643] = 8'h00;
reg_space[6644] = 8'h00;
reg_space[6645] = 8'h00;
reg_space[6646] = 8'h00;
reg_space[6647] = 8'h00;
reg_space[6648] = 8'h00;
reg_space[6649] = 8'h00;
reg_space[6650] = 8'h00;
reg_space[6651] = 8'h00;
reg_space[6652] = 8'h00;
reg_space[6653] = 8'h00;
reg_space[6654] = 8'h00;
reg_space[6655] = 8'h00;
reg_space[6656] = 8'h00;
reg_space[6657] = 8'h00;
reg_space[6658] = 8'h00;
reg_space[6659] = 8'h00;
reg_space[6660] = 8'h00;
reg_space[6661] = 8'h00;
reg_space[6662] = 8'h00;
reg_space[6663] = 8'h00;
reg_space[6664] = 8'h00;
reg_space[6665] = 8'h00;
reg_space[6666] = 8'h00;
reg_space[6667] = 8'h00;
reg_space[6668] = 8'h00;
reg_space[6669] = 8'h00;
reg_space[6670] = 8'h00;
reg_space[6671] = 8'h00;
reg_space[6672] = 8'h00;
reg_space[6673] = 8'h00;
reg_space[6674] = 8'h00;
reg_space[6675] = 8'h00;
reg_space[6676] = 8'h00;
reg_space[6677] = 8'h00;
reg_space[6678] = 8'h00;
reg_space[6679] = 8'h00;
reg_space[6680] = 8'h00;
reg_space[6681] = 8'h00;
reg_space[6682] = 8'h00;
reg_space[6683] = 8'h00;
reg_space[6684] = 8'h00;
reg_space[6685] = 8'h00;
reg_space[6686] = 8'h00;
reg_space[6687] = 8'h00;
reg_space[6688] = 8'h00;
reg_space[6689] = 8'h00;
reg_space[6690] = 8'h00;
reg_space[6691] = 8'h00;
reg_space[6692] = 8'h00;
reg_space[6693] = 8'h00;
reg_space[6694] = 8'h00;
reg_space[6695] = 8'h00;
reg_space[6696] = 8'h00;
reg_space[6697] = 8'h00;
reg_space[6698] = 8'h00;
reg_space[6699] = 8'h00;
reg_space[6700; = 8'h00;
reg_space[6701] = 8'h00;
reg_space[6702] = 8'h00;
reg_space[6703] = 8'h00;
reg_space[6704] = 8'h00;
reg_space[6705] = 8'h00;
reg_space[6706] = 8'h00;
reg_space[6707] = 8'h00;
reg_space[6708] = 8'h00;
reg_space[6709] = 8'h00;
reg_space[6710] = 8'h00;
reg_space[6711] = 8'h00;
reg_space[6712] = 8'h00;
reg_space[6713] = 8'h00;
reg_space[6714] = 8'h00;
reg_space[6715] = 8'h00;
reg_space[6716] = 8'h00;
reg_space[6717] = 8'h00;
reg_space[6718] = 8'h00;
reg_space[6719] = 8'h00;
reg_space[6720] = 8'h00;
reg_space[6721] = 8'h00;
reg_space[6722] = 8'h00;
reg_space[6723] = 8'h00;
reg_space[6724] = 8'h00;
reg_space[6725] = 8'h00;
reg_space[6726] = 8'h00;
reg_space[6727] = 8'h00;
reg_space[6728] = 8'h00;
reg_space[6729] = 8'h00;
reg_space[6730] = 8'h00;
reg_space[6731] = 8'h00;
reg_space[6732] = 8'h00;
reg_space[6733] = 8'h00;
reg_space[6734] = 8'h00;
reg_space[6735] = 8'h00;
reg_space[6736] = 8'h00;
reg_space[6737] = 8'h00;
reg_space[6738] = 8'h00;
reg_space[6739] = 8'h00;
reg_space[6740] = 8'h00;
reg_space[6741] = 8'h00;
reg_space[6742] = 8'h00;
reg_space[6743] = 8'h00;
reg_space[6744] = 8'h00;
reg_space[6745] = 8'h00;
reg_space[6746] = 8'h00;
reg_space[6747] = 8'h00;
reg_space[6748] = 8'h00;
reg_space[6749] = 8'h00;
reg_space[6750] = 8'h00;
reg_space[6751] = 8'h00;
reg_space[6752] = 8'h00;
reg_space[6753] = 8'h00;
reg_space[6754] = 8'h00;
reg_space[6755] = 8'h00;
reg_space[6756] = 8'h00;
reg_space[6757] = 8'h00;
reg_space[6758] = 8'h00;
reg_space[6759] = 8'h00;
reg_space[6760] = 8'h00;
reg_space[6761] = 8'h00;
reg_space[6762] = 8'h00;
reg_space[6763] = 8'h00;
reg_space[6764] = 8'h00;
reg_space[6765] = 8'h00;
reg_space[6766] = 8'h00;
reg_space[6767] = 8'h00;
reg_space[6768] = 8'h00;
reg_space[6769] = 8'h00;
reg_space[6770] = 8'h00;
reg_space[6771] = 8'h00;
reg_space[6772] = 8'h00;
reg_space[6773] = 8'h00;
reg_space[6774] = 8'h00;
reg_space[6775] = 8'h00;
reg_space[6776] = 8'h00;
reg_space[6777] = 8'h00;
reg_space[6778] = 8'h00;
reg_space[6779] = 8'h00;
reg_space[6780] = 8'h00;
reg_space[6781] = 8'h00;
reg_space[6782] = 8'h00;
reg_space[6783] = 8'h00;
reg_space[6784] = 8'h00;
reg_space[6785] = 8'h00;
reg_space[6786] = 8'h00;
reg_space[6787] = 8'h00;
reg_space[6788] = 8'h00;
reg_space[6789] = 8'h00;
reg_space[6790] = 8'h00;
reg_space[6791] = 8'h00;
reg_space[6792] = 8'h00;
reg_space[6793] = 8'h00;
reg_space[6794] = 8'h00;
reg_space[6795] = 8'h00;
reg_space[6796] = 8'h00;
reg_space[6797] = 8'h00;
reg_space[6798] = 8'h00;
reg_space[6799] = 8'h00;
reg_space[6800; = 8'h00;
reg_space[6801] = 8'h00;
reg_space[6802] = 8'h00;
reg_space[6803] = 8'h00;
reg_space[6804] = 8'h00;
reg_space[6805] = 8'h00;
reg_space[6806] = 8'h00;
reg_space[6807] = 8'h00;
reg_space[6808] = 8'h00;
reg_space[6809] = 8'h00;
reg_space[6810] = 8'h00;
reg_space[6811] = 8'h00;
reg_space[6812] = 8'h00;
reg_space[6813] = 8'h00;
reg_space[6814] = 8'h00;
reg_space[6815] = 8'h00;
reg_space[6816] = 8'h00;
reg_space[6817] = 8'h00;
reg_space[6818] = 8'h00;
reg_space[6819] = 8'h00;
reg_space[6820] = 8'h00;
reg_space[6821] = 8'h00;
reg_space[6822] = 8'h00;
reg_space[6823] = 8'h00;
reg_space[6824] = 8'h00;
reg_space[6825] = 8'h00;
reg_space[6826] = 8'h00;
reg_space[6827] = 8'h00;
reg_space[6828] = 8'h00;
reg_space[6829] = 8'h00;
reg_space[6830] = 8'h00;
reg_space[6831] = 8'h00;
reg_space[6832] = 8'h00;
reg_space[6833] = 8'h00;
reg_space[6834] = 8'h00;
reg_space[6835] = 8'h00;
reg_space[6836] = 8'h00;
reg_space[6837] = 8'h00;
reg_space[6838] = 8'h00;
reg_space[6839] = 8'h00;
reg_space[6840] = 8'h00;
reg_space[6841] = 8'h00;
reg_space[6842] = 8'h00;
reg_space[6843] = 8'h00;
reg_space[6844] = 8'h00;
reg_space[6845] = 8'h00;
reg_space[6846] = 8'h00;
reg_space[6847] = 8'h00;
reg_space[6848] = 8'h00;
reg_space[6849] = 8'h00;
reg_space[6850] = 8'h00;
reg_space[6851] = 8'h00;
reg_space[6852] = 8'h00;
reg_space[6853] = 8'h00;
reg_space[6854] = 8'h00;
reg_space[6855] = 8'h00;
reg_space[6856] = 8'h00;
reg_space[6857] = 8'h00;
reg_space[6858] = 8'h00;
reg_space[6859] = 8'h00;
reg_space[6860] = 8'h00;
reg_space[6861] = 8'h00;
reg_space[6862] = 8'h00;
reg_space[6863] = 8'h00;
reg_space[6864] = 8'h00;
reg_space[6865] = 8'h00;
reg_space[6866] = 8'h00;
reg_space[6867] = 8'h00;
reg_space[6868] = 8'h00;
reg_space[6869] = 8'h00;
reg_space[6870] = 8'h00;
reg_space[6871] = 8'h00;
reg_space[6872] = 8'h00;
reg_space[6873] = 8'h00;
reg_space[6874] = 8'h00;
reg_space[6875] = 8'h00;
reg_space[6876] = 8'h00;
reg_space[6877] = 8'h00;
reg_space[6878] = 8'h00;
reg_space[6879] = 8'h00;
reg_space[6880] = 8'h00;
reg_space[6881] = 8'h00;
reg_space[6882] = 8'h00;
reg_space[6883] = 8'h00;
reg_space[6884] = 8'h00;
reg_space[6885] = 8'h00;
reg_space[6886] = 8'h00;
reg_space[6887] = 8'h00;
reg_space[6888] = 8'h00;
reg_space[6889] = 8'h00;
reg_space[6890] = 8'h00;
reg_space[6891] = 8'h00;
reg_space[6892] = 8'h00;
reg_space[6893] = 8'h00;
reg_space[6894] = 8'h00;
reg_space[6895] = 8'h00;
reg_space[6896] = 8'h00;
reg_space[6897] = 8'h00;
reg_space[6898] = 8'h00;
reg_space[6899] = 8'h00;
reg_space[6900; = 8'h00;
reg_space[6901] = 8'h00;
reg_space[6902] = 8'h00;
reg_space[6903] = 8'h00;
reg_space[6904] = 8'h00;
reg_space[6905] = 8'h00;
reg_space[6906] = 8'h00;
reg_space[6907] = 8'h00;
reg_space[6908] = 8'h00;
reg_space[6909] = 8'h00;
reg_space[6910] = 8'h00;
reg_space[6911] = 8'h00;
reg_space[6912] = 8'h00;
reg_space[6913] = 8'h00;
reg_space[6914] = 8'h00;
reg_space[6915] = 8'h00;
reg_space[6916] = 8'h00;
reg_space[6917] = 8'h00;
reg_space[6918] = 8'h00;
reg_space[6919] = 8'h00;
reg_space[6920] = 8'h00;
reg_space[6921] = 8'h00;
reg_space[6922] = 8'h00;
reg_space[6923] = 8'h00;
reg_space[6924] = 8'h00;
reg_space[6925] = 8'h00;
reg_space[6926] = 8'h00;
reg_space[6927] = 8'h00;
reg_space[6928] = 8'h00;
reg_space[6929] = 8'h00;
reg_space[6930] = 8'h00;
reg_space[6931] = 8'h00;
reg_space[6932] = 8'h00;
reg_space[6933] = 8'h00;
reg_space[6934] = 8'h00;
reg_space[6935] = 8'h00;
reg_space[6936] = 8'h00;
reg_space[6937] = 8'h00;
reg_space[6938] = 8'h00;
reg_space[6939] = 8'h00;
reg_space[6940] = 8'h00;
reg_space[6941] = 8'h00;
reg_space[6942] = 8'h00;
reg_space[6943] = 8'h00;
reg_space[6944] = 8'h00;
reg_space[6945] = 8'h00;
reg_space[6946] = 8'h00;
reg_space[6947] = 8'h00;
reg_space[6948] = 8'h00;
reg_space[6949] = 8'h00;
reg_space[6950] = 8'h00;
reg_space[6951] = 8'h00;
reg_space[6952] = 8'h00;
reg_space[6953] = 8'h00;
reg_space[6954] = 8'h00;
reg_space[6955] = 8'h00;
reg_space[6956] = 8'h00;
reg_space[6957] = 8'h00;
reg_space[6958] = 8'h00;
reg_space[6959] = 8'h00;
reg_space[6960] = 8'h00;
reg_space[6961] = 8'h00;
reg_space[6962] = 8'h00;
reg_space[6963] = 8'h00;
reg_space[6964] = 8'h00;
reg_space[6965] = 8'h00;
reg_space[6966] = 8'h00;
reg_space[6967] = 8'h00;
reg_space[6968] = 8'h00;
reg_space[6969] = 8'h00;
reg_space[6970] = 8'h00;
reg_space[6971] = 8'h00;
reg_space[6972] = 8'h00;
reg_space[6973] = 8'h00;
reg_space[6974] = 8'h00;
reg_space[6975] = 8'h00;
reg_space[6976] = 8'h00;
reg_space[6977] = 8'h00;
reg_space[6978] = 8'h00;
reg_space[6979] = 8'h00;
reg_space[6980] = 8'h00;
reg_space[6981] = 8'h00;
reg_space[6982] = 8'h00;
reg_space[6983] = 8'h00;
reg_space[6984] = 8'h00;
reg_space[6985] = 8'h00;
reg_space[6986] = 8'h00;
reg_space[6987] = 8'h00;
reg_space[6988] = 8'h00;
reg_space[6989] = 8'h00;
reg_space[6990] = 8'h00;
reg_space[6991] = 8'h00;
reg_space[6992] = 8'h00;
reg_space[6993] = 8'h00;
reg_space[6994] = 8'h00;
reg_space[6995] = 8'h00;
reg_space[6996] = 8'h00;
reg_space[6997] = 8'h00;
reg_space[6998] = 8'h00;
reg_space[6999] = 8'h00;
reg_space[700;0] = 8'h00;
reg_space[700;1] = 8'h00;
reg_space[700;2] = 8'h00;
reg_space[700;3] = 8'h00;
reg_space[700;4] = 8'h00;
reg_space[700;5] = 8'h00;
reg_space[700;6] = 8'h00;
reg_space[700;7] = 8'h00;
reg_space[700;8] = 8'h00;
reg_space[700;9] = 8'h00;
reg_space[7010] = 8'h00;
reg_space[7011] = 8'h00;
reg_space[7012] = 8'h00;
reg_space[7013] = 8'h00;
reg_space[7014] = 8'h00;
reg_space[7015] = 8'h00;
reg_space[7016] = 8'h00;
reg_space[7017] = 8'h00;
reg_space[7018] = 8'h00;
reg_space[7019] = 8'h00;
reg_space[7020] = 8'h00;
reg_space[7021] = 8'h00;
reg_space[7022] = 8'h00;
reg_space[7023] = 8'h00;
reg_space[7024] = 8'h00;
reg_space[7025] = 8'h00;
reg_space[7026] = 8'h00;
reg_space[7027] = 8'h00;
reg_space[7028] = 8'h00;
reg_space[7029] = 8'h00;
reg_space[7030] = 8'h00;
reg_space[7031] = 8'h00;
reg_space[7032] = 8'h00;
reg_space[7033] = 8'h00;
reg_space[7034] = 8'h00;
reg_space[7035] = 8'h00;
reg_space[7036] = 8'h00;
reg_space[7037] = 8'h00;
reg_space[7038] = 8'h00;
reg_space[7039] = 8'h00;
reg_space[7040] = 8'h00;
reg_space[7041] = 8'h00;
reg_space[7042] = 8'h00;
reg_space[7043] = 8'h00;
reg_space[7044] = 8'h00;
reg_space[7045] = 8'h00;
reg_space[7046] = 8'h00;
reg_space[7047] = 8'h00;
reg_space[7048] = 8'h00;
reg_space[7049] = 8'h00;
reg_space[7050] = 8'h00;
reg_space[7051] = 8'h00;
reg_space[7052] = 8'h00;
reg_space[7053] = 8'h00;
reg_space[7054] = 8'h00;
reg_space[7055] = 8'h00;
reg_space[7056] = 8'h00;
reg_space[7057] = 8'h00;
reg_space[7058] = 8'h00;
reg_space[7059] = 8'h00;
reg_space[7060] = 8'h00;
reg_space[7061] = 8'h00;
reg_space[7062] = 8'h00;
reg_space[7063] = 8'h00;
reg_space[7064] = 8'h00;
reg_space[7065] = 8'h00;
reg_space[7066] = 8'h00;
reg_space[7067] = 8'h00;
reg_space[7068] = 8'h00;
reg_space[7069] = 8'h00;
reg_space[7070] = 8'h00;
reg_space[7071] = 8'h00;
reg_space[7072] = 8'h00;
reg_space[7073] = 8'h00;
reg_space[7074] = 8'h00;
reg_space[7075] = 8'h00;
reg_space[7076] = 8'h00;
reg_space[7077] = 8'h00;
reg_space[7078] = 8'h00;
reg_space[7079] = 8'h00;
reg_space[7080] = 8'h00;
reg_space[7081] = 8'h00;
reg_space[7082] = 8'h00;
reg_space[7083] = 8'h00;
reg_space[7084] = 8'h00;
reg_space[7085] = 8'h00;
reg_space[7086] = 8'h00;
reg_space[7087] = 8'h00;
reg_space[7088] = 8'h00;
reg_space[7089] = 8'h00;
reg_space[7090] = 8'h00;
reg_space[7091] = 8'h00;
reg_space[7092] = 8'h00;
reg_space[7093] = 8'h00;
reg_space[7094] = 8'h00;
reg_space[7095] = 8'h00;
reg_space[7096] = 8'h00;
reg_space[7097] = 8'h00;
reg_space[7098] = 8'h00;
reg_space[7099] = 8'h00;
reg_space[7100; = 8'h00;
reg_space[7101] = 8'h00;
reg_space[7102] = 8'h00;
reg_space[7103] = 8'h00;
reg_space[7104] = 8'h00;
reg_space[7105] = 8'h00;
reg_space[7106] = 8'h00;
reg_space[7107] = 8'h00;
reg_space[7108] = 8'h00;
reg_space[7109] = 8'h00;
reg_space[7110] = 8'h00;
reg_space[7111] = 8'h00;
reg_space[7112] = 8'h00;
reg_space[7113] = 8'h00;
reg_space[7114] = 8'h00;
reg_space[7115] = 8'h00;
reg_space[7116] = 8'h00;
reg_space[7117] = 8'h00;
reg_space[7118] = 8'h00;
reg_space[7119] = 8'h00;
reg_space[7120] = 8'h00;
reg_space[7121] = 8'h00;
reg_space[7122] = 8'h00;
reg_space[7123] = 8'h00;
reg_space[7124] = 8'h00;
reg_space[7125] = 8'h00;
reg_space[7126] = 8'h00;
reg_space[7127] = 8'h00;
reg_space[7128] = 8'h00;
reg_space[7129] = 8'h00;
reg_space[7130] = 8'h00;
reg_space[7131] = 8'h00;
reg_space[7132] = 8'h00;
reg_space[7133] = 8'h00;
reg_space[7134] = 8'h00;
reg_space[7135] = 8'h00;
reg_space[7136] = 8'h00;
reg_space[7137] = 8'h00;
reg_space[7138] = 8'h00;
reg_space[7139] = 8'h00;
reg_space[7140] = 8'h00;
reg_space[7141] = 8'h00;
reg_space[7142] = 8'h00;
reg_space[7143] = 8'h00;
reg_space[7144] = 8'h00;
reg_space[7145] = 8'h00;
reg_space[7146] = 8'h00;
reg_space[7147] = 8'h00;
reg_space[7148] = 8'h00;
reg_space[7149] = 8'h00;
reg_space[7150] = 8'h00;
reg_space[7151] = 8'h00;
reg_space[7152] = 8'h00;
reg_space[7153] = 8'h00;
reg_space[7154] = 8'h00;
reg_space[7155] = 8'h00;
reg_space[7156] = 8'h00;
reg_space[7157] = 8'h00;
reg_space[7158] = 8'h00;
reg_space[7159] = 8'h00;
reg_space[7160] = 8'h00;
reg_space[7161] = 8'h00;
reg_space[7162] = 8'h00;
reg_space[7163] = 8'h00;
reg_space[7164] = 8'h00;
reg_space[7165] = 8'h00;
reg_space[7166] = 8'h00;
reg_space[7167] = 8'h00;
reg_space[7168] = 8'h00;
reg_space[7169] = 8'h00;
reg_space[7170] = 8'h00;
reg_space[7171] = 8'h00;
reg_space[7172] = 8'h00;
reg_space[7173] = 8'h00;
reg_space[7174] = 8'h00;
reg_space[7175] = 8'h00;
reg_space[7176] = 8'h00;
reg_space[7177] = 8'h00;
reg_space[7178] = 8'h00;
reg_space[7179] = 8'h00;
reg_space[7180] = 8'h00;
reg_space[7181] = 8'h00;
reg_space[7182] = 8'h00;
reg_space[7183] = 8'h00;
reg_space[7184] = 8'h00;
reg_space[7185] = 8'h00;
reg_space[7186] = 8'h00;
reg_space[7187] = 8'h00;
reg_space[7188] = 8'h00;
reg_space[7189] = 8'h00;
reg_space[7190] = 8'h00;
reg_space[7191] = 8'h00;
reg_space[7192] = 8'h00;
reg_space[7193] = 8'h00;
reg_space[7194] = 8'h00;
reg_space[7195] = 8'h00;
reg_space[7196] = 8'h00;
reg_space[7197] = 8'h00;
reg_space[7198] = 8'h00;
reg_space[7199] = 8'h00;
reg_space[7200; = 8'h00;
reg_space[7201] = 8'h00;
reg_space[7202] = 8'h00;
reg_space[7203] = 8'h00;
reg_space[7204] = 8'h00;
reg_space[7205] = 8'h00;
reg_space[7206] = 8'h00;
reg_space[7207] = 8'h00;
reg_space[7208] = 8'h00;
reg_space[7209] = 8'h00;
reg_space[7210] = 8'h00;
reg_space[7211] = 8'h00;
reg_space[7212] = 8'h00;
reg_space[7213] = 8'h00;
reg_space[7214] = 8'h00;
reg_space[7215] = 8'h00;
reg_space[7216] = 8'h00;
reg_space[7217] = 8'h00;
reg_space[7218] = 8'h00;
reg_space[7219] = 8'h00;
reg_space[7220] = 8'h00;
reg_space[7221] = 8'h00;
reg_space[7222] = 8'h00;
reg_space[7223] = 8'h00;
reg_space[7224] = 8'h00;
reg_space[7225] = 8'h00;
reg_space[7226] = 8'h00;
reg_space[7227] = 8'h00;
reg_space[7228] = 8'h00;
reg_space[7229] = 8'h00;
reg_space[7230] = 8'h00;
reg_space[7231] = 8'h00;
reg_space[7232] = 8'h00;
reg_space[7233] = 8'h00;
reg_space[7234] = 8'h00;
reg_space[7235] = 8'h00;
reg_space[7236] = 8'h00;
reg_space[7237] = 8'h00;
reg_space[7238] = 8'h00;
reg_space[7239] = 8'h00;
reg_space[7240] = 8'h00;
reg_space[7241] = 8'h00;
reg_space[7242] = 8'h00;
reg_space[7243] = 8'h00;
reg_space[7244] = 8'h00;
reg_space[7245] = 8'h00;
reg_space[7246] = 8'h00;
reg_space[7247] = 8'h00;
reg_space[7248] = 8'h00;
reg_space[7249] = 8'h00;
reg_space[7250] = 8'h00;
reg_space[7251] = 8'h00;
reg_space[7252] = 8'h00;
reg_space[7253] = 8'h00;
reg_space[7254] = 8'h00;
reg_space[7255] = 8'h00;
reg_space[7256] = 8'h00;
reg_space[7257] = 8'h00;
reg_space[7258] = 8'h00;
reg_space[7259] = 8'h00;
reg_space[7260] = 8'h00;
reg_space[7261] = 8'h00;
reg_space[7262] = 8'h00;
reg_space[7263] = 8'h00;
reg_space[7264] = 8'h00;
reg_space[7265] = 8'h00;
reg_space[7266] = 8'h00;
reg_space[7267] = 8'h00;
reg_space[7268] = 8'h00;
reg_space[7269] = 8'h00;
reg_space[7270] = 8'h00;
reg_space[7271] = 8'h00;
reg_space[7272] = 8'h00;
reg_space[7273] = 8'h00;
reg_space[7274] = 8'h00;
reg_space[7275] = 8'h00;
reg_space[7276] = 8'h00;
reg_space[7277] = 8'h00;
reg_space[7278] = 8'h00;
reg_space[7279] = 8'h00;
reg_space[7280] = 8'h00;
reg_space[7281] = 8'h00;
reg_space[7282] = 8'h00;
reg_space[7283] = 8'h00;
reg_space[7284] = 8'h00;
reg_space[7285] = 8'h00;
reg_space[7286] = 8'h00;
reg_space[7287] = 8'h00;
reg_space[7288] = 8'h00;
reg_space[7289] = 8'h00;
reg_space[7290] = 8'h00;
reg_space[7291] = 8'h00;
reg_space[7292] = 8'h00;
reg_space[7293] = 8'h00;
reg_space[7294] = 8'h00;
reg_space[7295] = 8'h00;
reg_space[7296] = 8'h00;
reg_space[7297] = 8'h00;
reg_space[7298] = 8'h00;
reg_space[7299] = 8'h00;
reg_space[7300; = 8'h00;
reg_space[7301] = 8'h00;
reg_space[7302] = 8'h00;
reg_space[7303] = 8'h00;
reg_space[7304] = 8'h00;
reg_space[7305] = 8'h00;
reg_space[7306] = 8'h00;
reg_space[7307] = 8'h00;
reg_space[7308] = 8'h00;
reg_space[7309] = 8'h00;
reg_space[7310] = 8'h00;
reg_space[7311] = 8'h00;
reg_space[7312] = 8'h00;
reg_space[7313] = 8'h00;
reg_space[7314] = 8'h00;
reg_space[7315] = 8'h00;
reg_space[7316] = 8'h00;
reg_space[7317] = 8'h00;
reg_space[7318] = 8'h00;
reg_space[7319] = 8'h00;
reg_space[7320] = 8'h00;
reg_space[7321] = 8'h00;
reg_space[7322] = 8'h00;
reg_space[7323] = 8'h00;
reg_space[7324] = 8'h00;
reg_space[7325] = 8'h00;
reg_space[7326] = 8'h00;
reg_space[7327] = 8'h00;
reg_space[7328] = 8'h00;
reg_space[7329] = 8'h00;
reg_space[7330] = 8'h00;
reg_space[7331] = 8'h00;
reg_space[7332] = 8'h00;
reg_space[7333] = 8'h00;
reg_space[7334] = 8'h00;
reg_space[7335] = 8'h00;
reg_space[7336] = 8'h00;
reg_space[7337] = 8'h00;
reg_space[7338] = 8'h00;
reg_space[7339] = 8'h00;
reg_space[7340] = 8'h00;
reg_space[7341] = 8'h00;
reg_space[7342] = 8'h00;
reg_space[7343] = 8'h00;
reg_space[7344] = 8'h00;
reg_space[7345] = 8'h00;
reg_space[7346] = 8'h00;
reg_space[7347] = 8'h00;
reg_space[7348] = 8'h00;
reg_space[7349] = 8'h00;
reg_space[7350] = 8'h00;
reg_space[7351] = 8'h00;
reg_space[7352] = 8'h00;
reg_space[7353] = 8'h00;
reg_space[7354] = 8'h00;
reg_space[7355] = 8'h00;
reg_space[7356] = 8'h00;
reg_space[7357] = 8'h00;
reg_space[7358] = 8'h00;
reg_space[7359] = 8'h00;
reg_space[7360] = 8'h00;
reg_space[7361] = 8'h00;
reg_space[7362] = 8'h00;
reg_space[7363] = 8'h00;
reg_space[7364] = 8'h00;
reg_space[7365] = 8'h00;
reg_space[7366] = 8'h00;
reg_space[7367] = 8'h00;
reg_space[7368] = 8'h00;
reg_space[7369] = 8'h00;
reg_space[7370] = 8'h00;
reg_space[7371] = 8'h00;
reg_space[7372] = 8'h00;
reg_space[7373] = 8'h00;
reg_space[7374] = 8'h00;
reg_space[7375] = 8'h00;
reg_space[7376] = 8'h00;
reg_space[7377] = 8'h00;
reg_space[7378] = 8'h00;
reg_space[7379] = 8'h00;
reg_space[7380] = 8'h00;
reg_space[7381] = 8'h00;
reg_space[7382] = 8'h00;
reg_space[7383] = 8'h00;
reg_space[7384] = 8'h00;
reg_space[7385] = 8'h00;
reg_space[7386] = 8'h00;
reg_space[7387] = 8'h00;
reg_space[7388] = 8'h00;
reg_space[7389] = 8'h00;
reg_space[7390] = 8'h00;
reg_space[7391] = 8'h00;
reg_space[7392] = 8'h00;
reg_space[7393] = 8'h00;
reg_space[7394] = 8'h00;
reg_space[7395] = 8'h00;
reg_space[7396] = 8'h00;
reg_space[7397] = 8'h00;
reg_space[7398] = 8'h00;
reg_space[7399] = 8'h00;
reg_space[7400; = 8'h00;
reg_space[7401] = 8'h00;
reg_space[7402] = 8'h00;
reg_space[7403] = 8'h00;
reg_space[7404] = 8'h00;
reg_space[7405] = 8'h00;
reg_space[7406] = 8'h00;
reg_space[7407] = 8'h00;
reg_space[7408] = 8'h00;
reg_space[7409] = 8'h00;
reg_space[7410] = 8'h00;
reg_space[7411] = 8'h00;
reg_space[7412] = 8'h00;
reg_space[7413] = 8'h00;
reg_space[7414] = 8'h00;
reg_space[7415] = 8'h00;
reg_space[7416] = 8'h00;
reg_space[7417] = 8'h00;
reg_space[7418] = 8'h00;
reg_space[7419] = 8'h00;
reg_space[7420] = 8'h00;
reg_space[7421] = 8'h00;
reg_space[7422] = 8'h00;
reg_space[7423] = 8'h00;
reg_space[7424] = 8'h00;
reg_space[7425] = 8'h00;
reg_space[7426] = 8'h00;
reg_space[7427] = 8'h00;
reg_space[7428] = 8'h00;
reg_space[7429] = 8'h00;
reg_space[7430] = 8'h00;
reg_space[7431] = 8'h00;
reg_space[7432] = 8'h00;
reg_space[7433] = 8'h00;
reg_space[7434] = 8'h00;
reg_space[7435] = 8'h00;
reg_space[7436] = 8'h00;
reg_space[7437] = 8'h00;
reg_space[7438] = 8'h00;
reg_space[7439] = 8'h00;
reg_space[7440] = 8'h00;
reg_space[7441] = 8'h00;
reg_space[7442] = 8'h00;
reg_space[7443] = 8'h00;
reg_space[7444] = 8'h00;
reg_space[7445] = 8'h00;
reg_space[7446] = 8'h00;
reg_space[7447] = 8'h00;
reg_space[7448] = 8'h00;
reg_space[7449] = 8'h00;
reg_space[7450] = 8'h00;
reg_space[7451] = 8'h00;
reg_space[7452] = 8'h00;
reg_space[7453] = 8'h00;
reg_space[7454] = 8'h00;
reg_space[7455] = 8'h00;
reg_space[7456] = 8'h00;
reg_space[7457] = 8'h00;
reg_space[7458] = 8'h00;
reg_space[7459] = 8'h00;
reg_space[7460] = 8'h00;
reg_space[7461] = 8'h00;
reg_space[7462] = 8'h00;
reg_space[7463] = 8'h00;
reg_space[7464] = 8'h00;
reg_space[7465] = 8'h00;
reg_space[7466] = 8'h00;
reg_space[7467] = 8'h00;
reg_space[7468] = 8'h00;
reg_space[7469] = 8'h00;
reg_space[7470] = 8'h00;
reg_space[7471] = 8'h00;
reg_space[7472] = 8'h00;
reg_space[7473] = 8'h00;
reg_space[7474] = 8'h00;
reg_space[7475] = 8'h00;
reg_space[7476] = 8'h00;
reg_space[7477] = 8'h00;
reg_space[7478] = 8'h00;
reg_space[7479] = 8'h00;
reg_space[7480] = 8'h00;
reg_space[7481] = 8'h00;
reg_space[7482] = 8'h00;
reg_space[7483] = 8'h00;
reg_space[7484] = 8'h00;
reg_space[7485] = 8'h00;
reg_space[7486] = 8'h00;
reg_space[7487] = 8'h00;
reg_space[7488] = 8'h00;
reg_space[7489] = 8'h00;
reg_space[7490] = 8'h00;
reg_space[7491] = 8'h00;
reg_space[7492] = 8'h00;
reg_space[7493] = 8'h00;
reg_space[7494] = 8'h00;
reg_space[7495] = 8'h00;
reg_space[7496] = 8'h00;
reg_space[7497] = 8'h00;
reg_space[7498] = 8'h00;
reg_space[7499] = 8'h00;
reg_space[7500; = 8'h00;
reg_space[7501] = 8'h00;
reg_space[7502] = 8'h00;
reg_space[7503] = 8'h00;
reg_space[7504] = 8'h00;
reg_space[7505] = 8'h00;
reg_space[7506] = 8'h00;
reg_space[7507] = 8'h00;
reg_space[7508] = 8'h00;
reg_space[7509] = 8'h00;
reg_space[7510] = 8'h00;
reg_space[7511] = 8'h00;
reg_space[7512] = 8'h00;
reg_space[7513] = 8'h00;
reg_space[7514] = 8'h00;
reg_space[7515] = 8'h00;
reg_space[7516] = 8'h00;
reg_space[7517] = 8'h00;
reg_space[7518] = 8'h00;
reg_space[7519] = 8'h00;
reg_space[7520] = 8'h00;
reg_space[7521] = 8'h00;
reg_space[7522] = 8'h00;
reg_space[7523] = 8'h00;
reg_space[7524] = 8'h00;
reg_space[7525] = 8'h00;
reg_space[7526] = 8'h00;
reg_space[7527] = 8'h00;
reg_space[7528] = 8'h00;
reg_space[7529] = 8'h00;
reg_space[7530] = 8'h00;
reg_space[7531] = 8'h00;
reg_space[7532] = 8'h00;
reg_space[7533] = 8'h00;
reg_space[7534] = 8'h00;
reg_space[7535] = 8'h00;
reg_space[7536] = 8'h00;
reg_space[7537] = 8'h00;
reg_space[7538] = 8'h00;
reg_space[7539] = 8'h00;
reg_space[7540] = 8'h00;
reg_space[7541] = 8'h00;
reg_space[7542] = 8'h00;
reg_space[7543] = 8'h00;
reg_space[7544] = 8'h00;
reg_space[7545] = 8'h00;
reg_space[7546] = 8'h00;
reg_space[7547] = 8'h00;
reg_space[7548] = 8'h00;
reg_space[7549] = 8'h00;
reg_space[7550] = 8'h00;
reg_space[7551] = 8'h00;
reg_space[7552] = 8'h00;
reg_space[7553] = 8'h00;
reg_space[7554] = 8'h00;
reg_space[7555] = 8'h00;
reg_space[7556] = 8'h00;
reg_space[7557] = 8'h00;
reg_space[7558] = 8'h00;
reg_space[7559] = 8'h00;
reg_space[7560] = 8'h00;
reg_space[7561] = 8'h00;
reg_space[7562] = 8'h00;
reg_space[7563] = 8'h00;
reg_space[7564] = 8'h00;
reg_space[7565] = 8'h00;
reg_space[7566] = 8'h00;
reg_space[7567] = 8'h00;
reg_space[7568] = 8'h00;
reg_space[7569] = 8'h00;
reg_space[7570] = 8'h00;
reg_space[7571] = 8'h00;
reg_space[7572] = 8'h00;
reg_space[7573] = 8'h00;
reg_space[7574] = 8'h00;
reg_space[7575] = 8'h00;
reg_space[7576] = 8'h00;
reg_space[7577] = 8'h00;
reg_space[7578] = 8'h00;
reg_space[7579] = 8'h00;
reg_space[7580] = 8'h00;
reg_space[7581] = 8'h00;
reg_space[7582] = 8'h00;
reg_space[7583] = 8'h00;
reg_space[7584] = 8'h00;
reg_space[7585] = 8'h00;
reg_space[7586] = 8'h00;
reg_space[7587] = 8'h00;
reg_space[7588] = 8'h00;
reg_space[7589] = 8'h00;
reg_space[7590] = 8'h00;
reg_space[7591] = 8'h00;
reg_space[7592] = 8'h00;
reg_space[7593] = 8'h00;
reg_space[7594] = 8'h00;
reg_space[7595] = 8'h00;
reg_space[7596] = 8'h00;
reg_space[7597] = 8'h00;
reg_space[7598] = 8'h00;
reg_space[7599] = 8'h00;
reg_space[7600; = 8'h00;
reg_space[7601] = 8'h00;
reg_space[7602] = 8'h00;
reg_space[7603] = 8'h00;
reg_space[7604] = 8'h00;
reg_space[7605] = 8'h00;
reg_space[7606] = 8'h00;
reg_space[7607] = 8'h00;
reg_space[7608] = 8'h00;
reg_space[7609] = 8'h00;
reg_space[7610] = 8'h00;
reg_space[7611] = 8'h00;
reg_space[7612] = 8'h00;
reg_space[7613] = 8'h00;
reg_space[7614] = 8'h00;
reg_space[7615] = 8'h00;
reg_space[7616] = 8'h00;
reg_space[7617] = 8'h00;
reg_space[7618] = 8'h00;
reg_space[7619] = 8'h00;
reg_space[7620] = 8'h00;
reg_space[7621] = 8'h00;
reg_space[7622] = 8'h00;
reg_space[7623] = 8'h00;
reg_space[7624] = 8'h00;
reg_space[7625] = 8'h00;
reg_space[7626] = 8'h00;
reg_space[7627] = 8'h00;
reg_space[7628] = 8'h00;
reg_space[7629] = 8'h00;
reg_space[7630] = 8'h00;
reg_space[7631] = 8'h00;
reg_space[7632] = 8'h00;
reg_space[7633] = 8'h00;
reg_space[7634] = 8'h00;
reg_space[7635] = 8'h00;
reg_space[7636] = 8'h00;
reg_space[7637] = 8'h00;
reg_space[7638] = 8'h00;
reg_space[7639] = 8'h00;
reg_space[7640] = 8'h00;
reg_space[7641] = 8'h00;
reg_space[7642] = 8'h00;
reg_space[7643] = 8'h00;
reg_space[7644] = 8'h00;
reg_space[7645] = 8'h00;
reg_space[7646] = 8'h00;
reg_space[7647] = 8'h00;
reg_space[7648] = 8'h00;
reg_space[7649] = 8'h00;
reg_space[7650] = 8'h00;
reg_space[7651] = 8'h00;
reg_space[7652] = 8'h00;
reg_space[7653] = 8'h00;
reg_space[7654] = 8'h00;
reg_space[7655] = 8'h00;
reg_space[7656] = 8'h00;
reg_space[7657] = 8'h00;
reg_space[7658] = 8'h00;
reg_space[7659] = 8'h00;
reg_space[7660] = 8'h00;
reg_space[7661] = 8'h00;
reg_space[7662] = 8'h00;
reg_space[7663] = 8'h00;
reg_space[7664] = 8'h00;
reg_space[7665] = 8'h00;
reg_space[7666] = 8'h00;
reg_space[7667] = 8'h00;
reg_space[7668] = 8'h00;
reg_space[7669] = 8'h00;
reg_space[7670] = 8'h00;
reg_space[7671] = 8'h00;
reg_space[7672] = 8'h00;
reg_space[7673] = 8'h00;
reg_space[7674] = 8'h00;
reg_space[7675] = 8'h00;
reg_space[7676] = 8'h00;
reg_space[7677] = 8'h00;
reg_space[7678] = 8'h00;
reg_space[7679] = 8'h00;
reg_space[7680] = 8'h00;
reg_space[7681] = 8'h00;
reg_space[7682] = 8'h00;
reg_space[7683] = 8'h00;
reg_space[7684] = 8'h00;
reg_space[7685] = 8'h00;
reg_space[7686] = 8'h00;
reg_space[7687] = 8'h00;
reg_space[7688] = 8'h00;
reg_space[7689] = 8'h00;
reg_space[7690] = 8'h00;
reg_space[7691] = 8'h00;
reg_space[7692] = 8'h00;
reg_space[7693] = 8'h00;
reg_space[7694] = 8'h00;
reg_space[7695] = 8'h00;
reg_space[7696] = 8'h00;
reg_space[7697] = 8'h00;
reg_space[7698] = 8'h00;
reg_space[7699] = 8'h00;
reg_space[7700; = 8'h00;
reg_space[7701] = 8'h00;
reg_space[7702] = 8'h00;
reg_space[7703] = 8'h00;
reg_space[7704] = 8'h00;
reg_space[7705] = 8'h00;
reg_space[7706] = 8'h00;
reg_space[7707] = 8'h00;
reg_space[7708] = 8'h00;
reg_space[7709] = 8'h00;
reg_space[7710] = 8'h00;
reg_space[7711] = 8'h00;
reg_space[7712] = 8'h00;
reg_space[7713] = 8'h00;
reg_space[7714] = 8'h00;
reg_space[7715] = 8'h00;
reg_space[7716] = 8'h00;
reg_space[7717] = 8'h00;
reg_space[7718] = 8'h00;
reg_space[7719] = 8'h00;
reg_space[7720] = 8'h00;
reg_space[7721] = 8'h00;
reg_space[7722] = 8'h00;
reg_space[7723] = 8'h00;
reg_space[7724] = 8'h00;
reg_space[7725] = 8'h00;
reg_space[7726] = 8'h00;
reg_space[7727] = 8'h00;
reg_space[7728] = 8'h00;
reg_space[7729] = 8'h00;
reg_space[7730] = 8'h00;
reg_space[7731] = 8'h00;
reg_space[7732] = 8'h00;
reg_space[7733] = 8'h00;
reg_space[7734] = 8'h00;
reg_space[7735] = 8'h00;
reg_space[7736] = 8'h00;
reg_space[7737] = 8'h00;
reg_space[7738] = 8'h00;
reg_space[7739] = 8'h00;
reg_space[7740] = 8'h00;
reg_space[7741] = 8'h00;
reg_space[7742] = 8'h00;
reg_space[7743] = 8'h00;
reg_space[7744] = 8'h00;
reg_space[7745] = 8'h00;
reg_space[7746] = 8'h00;
reg_space[7747] = 8'h00;
reg_space[7748] = 8'h00;
reg_space[7749] = 8'h00;
reg_space[7750] = 8'h00;
reg_space[7751] = 8'h00;
reg_space[7752] = 8'h00;
reg_space[7753] = 8'h00;
reg_space[7754] = 8'h00;
reg_space[7755] = 8'h00;
reg_space[7756] = 8'h00;
reg_space[7757] = 8'h00;
reg_space[7758] = 8'h00;
reg_space[7759] = 8'h00;
reg_space[7760] = 8'h00;
reg_space[7761] = 8'h00;
reg_space[7762] = 8'h00;
reg_space[7763] = 8'h00;
reg_space[7764] = 8'h00;
reg_space[7765] = 8'h00;
reg_space[7766] = 8'h00;
reg_space[7767] = 8'h00;
reg_space[7768] = 8'h00;
reg_space[7769] = 8'h00;
reg_space[7770] = 8'h00;
reg_space[7771] = 8'h00;
reg_space[7772] = 8'h00;
reg_space[7773] = 8'h00;
reg_space[7774] = 8'h00;
reg_space[7775] = 8'h00;
reg_space[7776] = 8'h00;
reg_space[7777] = 8'h00;
reg_space[7778] = 8'h00;
reg_space[7779] = 8'h00;
reg_space[7780] = 8'h00;
reg_space[7781] = 8'h00;
reg_space[7782] = 8'h00;
reg_space[7783] = 8'h00;
reg_space[7784] = 8'h00;
reg_space[7785] = 8'h00;
reg_space[7786] = 8'h00;
reg_space[7787] = 8'h00;
reg_space[7788] = 8'h00;
reg_space[7789] = 8'h00;
reg_space[7790] = 8'h00;
reg_space[7791] = 8'h00;
reg_space[7792] = 8'h00;
reg_space[7793] = 8'h00;
reg_space[7794] = 8'h00;
reg_space[7795] = 8'h00;
reg_space[7796] = 8'h00;
reg_space[7797] = 8'h00;
reg_space[7798] = 8'h00;
reg_space[7799] = 8'h00;
reg_space[7800; = 8'h00;
reg_space[7801] = 8'h00;
reg_space[7802] = 8'h00;
reg_space[7803] = 8'h00;
reg_space[7804] = 8'h00;
reg_space[7805] = 8'h00;
reg_space[7806] = 8'h00;
reg_space[7807] = 8'h00;
reg_space[7808] = 8'h00;
reg_space[7809] = 8'h00;
reg_space[7810] = 8'h00;
reg_space[7811] = 8'h00;
reg_space[7812] = 8'h00;
reg_space[7813] = 8'h00;
reg_space[7814] = 8'h00;
reg_space[7815] = 8'h00;
reg_space[7816] = 8'h00;
reg_space[7817] = 8'h00;
reg_space[7818] = 8'h00;
reg_space[7819] = 8'h00;
reg_space[7820] = 8'h00;
reg_space[7821] = 8'h00;
reg_space[7822] = 8'h00;
reg_space[7823] = 8'h00;
reg_space[7824] = 8'h00;
reg_space[7825] = 8'h00;
reg_space[7826] = 8'h00;
reg_space[7827] = 8'h00;
reg_space[7828] = 8'h00;
reg_space[7829] = 8'h00;
reg_space[7830] = 8'h00;
reg_space[7831] = 8'h00;
reg_space[7832] = 8'h00;
reg_space[7833] = 8'h00;
reg_space[7834] = 8'h00;
reg_space[7835] = 8'h00;
reg_space[7836] = 8'h00;
reg_space[7837] = 8'h00;
reg_space[7838] = 8'h00;
reg_space[7839] = 8'h00;
reg_space[7840] = 8'h00;
reg_space[7841] = 8'h00;
reg_space[7842] = 8'h00;
reg_space[7843] = 8'h00;
reg_space[7844] = 8'h00;
reg_space[7845] = 8'h00;
reg_space[7846] = 8'h00;
reg_space[7847] = 8'h00;
reg_space[7848] = 8'h00;
reg_space[7849] = 8'h00;
reg_space[7850] = 8'h00;
reg_space[7851] = 8'h00;
reg_space[7852] = 8'h00;
reg_space[7853] = 8'h00;
reg_space[7854] = 8'h00;
reg_space[7855] = 8'h00;
reg_space[7856] = 8'h00;
reg_space[7857] = 8'h00;
reg_space[7858] = 8'h00;
reg_space[7859] = 8'h00;
reg_space[7860] = 8'h00;
reg_space[7861] = 8'h00;
reg_space[7862] = 8'h00;
reg_space[7863] = 8'h00;
reg_space[7864] = 8'h00;
reg_space[7865] = 8'h00;
reg_space[7866] = 8'h00;
reg_space[7867] = 8'h00;
reg_space[7868] = 8'h00;
reg_space[7869] = 8'h00;
reg_space[7870] = 8'h00;
reg_space[7871] = 8'h00;
reg_space[7872] = 8'h00;
reg_space[7873] = 8'h00;
reg_space[7874] = 8'h00;
reg_space[7875] = 8'h00;
reg_space[7876] = 8'h00;
reg_space[7877] = 8'h00;
reg_space[7878] = 8'h00;
reg_space[7879] = 8'h00;
reg_space[7880] = 8'h00;
reg_space[7881] = 8'h00;
reg_space[7882] = 8'h00;
reg_space[7883] = 8'h00;
reg_space[7884] = 8'h00;
reg_space[7885] = 8'h00;
reg_space[7886] = 8'h00;
reg_space[7887] = 8'h00;
reg_space[7888] = 8'h00;
reg_space[7889] = 8'h00;
reg_space[7890] = 8'h00;
reg_space[7891] = 8'h00;
reg_space[7892] = 8'h00;
reg_space[7893] = 8'h00;
reg_space[7894] = 8'h00;
reg_space[7895] = 8'h00;
reg_space[7896] = 8'h00;
reg_space[7897] = 8'h00;
reg_space[7898] = 8'h00;
reg_space[7899] = 8'h00;
reg_space[7900; = 8'h00;
reg_space[7901] = 8'h00;
reg_space[7902] = 8'h00;
reg_space[7903] = 8'h00;
reg_space[7904] = 8'h00;
reg_space[7905] = 8'h00;
reg_space[7906] = 8'h00;
reg_space[7907] = 8'h00;
reg_space[7908] = 8'h00;
reg_space[7909] = 8'h00;
reg_space[7910] = 8'h00;
reg_space[7911] = 8'h00;
reg_space[7912] = 8'h00;
reg_space[7913] = 8'h00;
reg_space[7914] = 8'h00;
reg_space[7915] = 8'h00;
reg_space[7916] = 8'h00;
reg_space[7917] = 8'h00;
reg_space[7918] = 8'h00;
reg_space[7919] = 8'h00;
reg_space[7920] = 8'h00;
reg_space[7921] = 8'h00;
reg_space[7922] = 8'h00;
reg_space[7923] = 8'h00;
reg_space[7924] = 8'h00;
reg_space[7925] = 8'h00;
reg_space[7926] = 8'h00;
reg_space[7927] = 8'h00;
reg_space[7928] = 8'h00;
reg_space[7929] = 8'h00;
reg_space[7930] = 8'h00;
reg_space[7931] = 8'h00;
reg_space[7932] = 8'h00;
reg_space[7933] = 8'h00;
reg_space[7934] = 8'h00;
reg_space[7935] = 8'h00;
reg_space[7936] = 8'h00;
reg_space[7937] = 8'h00;
reg_space[7938] = 8'h00;
reg_space[7939] = 8'h00;
reg_space[7940] = 8'h00;
reg_space[7941] = 8'h00;
reg_space[7942] = 8'h00;
reg_space[7943] = 8'h00;
reg_space[7944] = 8'h00;
reg_space[7945] = 8'h00;
reg_space[7946] = 8'h00;
reg_space[7947] = 8'h00;
reg_space[7948] = 8'h00;
reg_space[7949] = 8'h00;
reg_space[7950] = 8'h00;
reg_space[7951] = 8'h00;
reg_space[7952] = 8'h00;
reg_space[7953] = 8'h00;
reg_space[7954] = 8'h00;
reg_space[7955] = 8'h00;
reg_space[7956] = 8'h00;
reg_space[7957] = 8'h00;
reg_space[7958] = 8'h00;
reg_space[7959] = 8'h00;
reg_space[7960] = 8'h00;
reg_space[7961] = 8'h00;
reg_space[7962] = 8'h00;
reg_space[7963] = 8'h00;
reg_space[7964] = 8'h00;
reg_space[7965] = 8'h00;
reg_space[7966] = 8'h00;
reg_space[7967] = 8'h00;
reg_space[7968] = 8'h00;
reg_space[7969] = 8'h00;
reg_space[7970] = 8'h00;
reg_space[7971] = 8'h00;
reg_space[7972] = 8'h00;
reg_space[7973] = 8'h00;
reg_space[7974] = 8'h00;
reg_space[7975] = 8'h00;
reg_space[7976] = 8'h00;
reg_space[7977] = 8'h00;
reg_space[7978] = 8'h00;
reg_space[7979] = 8'h00;
reg_space[7980] = 8'h00;
reg_space[7981] = 8'h00;
reg_space[7982] = 8'h00;
reg_space[7983] = 8'h00;
reg_space[7984] = 8'h00;
reg_space[7985] = 8'h00;
reg_space[7986] = 8'h00;
reg_space[7987] = 8'h00;
reg_space[7988] = 8'h00;
reg_space[7989] = 8'h00;
reg_space[7990] = 8'h00;
reg_space[7991] = 8'h00;
reg_space[7992] = 8'h00;
reg_space[7993] = 8'h00;
reg_space[7994] = 8'h00;
reg_space[7995] = 8'h00;
reg_space[7996] = 8'h00;
reg_space[7997] = 8'h00;
reg_space[7998] = 8'h00;
reg_space[7999] = 8'h00;
reg_space[800;0] = 8'h00;
reg_space[800;1] = 8'h00;
reg_space[800;2] = 8'h00;
reg_space[800;3] = 8'h00;
reg_space[800;4] = 8'h00;
reg_space[800;5] = 8'h00;
reg_space[800;6] = 8'h00;
reg_space[800;7] = 8'h00;
reg_space[800;8] = 8'h00;
reg_space[800;9] = 8'h00;
reg_space[8010] = 8'h00;
reg_space[8011] = 8'h00;
reg_space[8012] = 8'h00;
reg_space[8013] = 8'h00;
reg_space[8014] = 8'h00;
reg_space[8015] = 8'h00;
reg_space[8016] = 8'h00;
reg_space[8017] = 8'h00;
reg_space[8018] = 8'h00;
reg_space[8019] = 8'h00;
reg_space[8020] = 8'h00;
reg_space[8021] = 8'h00;
reg_space[8022] = 8'h00;
reg_space[8023] = 8'h00;
reg_space[8024] = 8'h00;
reg_space[8025] = 8'h00;
reg_space[8026] = 8'h00;
reg_space[8027] = 8'h00;
reg_space[8028] = 8'h00;
reg_space[8029] = 8'h00;
reg_space[8030] = 8'h00;
reg_space[8031] = 8'h00;
reg_space[8032] = 8'h00;
reg_space[8033] = 8'h00;
reg_space[8034] = 8'h00;
reg_space[8035] = 8'h00;
reg_space[8036] = 8'h00;
reg_space[8037] = 8'h00;
reg_space[8038] = 8'h00;
reg_space[8039] = 8'h00;
reg_space[8040] = 8'h00;
reg_space[8041] = 8'h00;
reg_space[8042] = 8'h00;
reg_space[8043] = 8'h00;
reg_space[8044] = 8'h00;
reg_space[8045] = 8'h00;
reg_space[8046] = 8'h00;
reg_space[8047] = 8'h00;
reg_space[8048] = 8'h00;
reg_space[8049] = 8'h00;
reg_space[8050] = 8'h00;
reg_space[8051] = 8'h00;
reg_space[8052] = 8'h00;
reg_space[8053] = 8'h00;
reg_space[8054] = 8'h00;
reg_space[8055] = 8'h00;
reg_space[8056] = 8'h00;
reg_space[8057] = 8'h00;
reg_space[8058] = 8'h00;
reg_space[8059] = 8'h00;
reg_space[8060] = 8'h00;
reg_space[8061] = 8'h00;
reg_space[8062] = 8'h00;
reg_space[8063] = 8'h00;
reg_space[8064] = 8'h00;
reg_space[8065] = 8'h00;
reg_space[8066] = 8'h00;
reg_space[8067] = 8'h00;
reg_space[8068] = 8'h00;
reg_space[8069] = 8'h00;
reg_space[8070] = 8'h00;
reg_space[8071] = 8'h00;
reg_space[8072] = 8'h00;
reg_space[8073] = 8'h00;
reg_space[8074] = 8'h00;
reg_space[8075] = 8'h00;
reg_space[8076] = 8'h00;
reg_space[8077] = 8'h00;
reg_space[8078] = 8'h00;
reg_space[8079] = 8'h00;
reg_space[8080] = 8'h00;
reg_space[8081] = 8'h00;
reg_space[8082] = 8'h00;
reg_space[8083] = 8'h00;
reg_space[8084] = 8'h00;
reg_space[8085] = 8'h00;
reg_space[8086] = 8'h00;
reg_space[8087] = 8'h00;
reg_space[8088] = 8'h00;
reg_space[8089] = 8'h00;
reg_space[8090] = 8'h00;
reg_space[8091] = 8'h00;
reg_space[8092] = 8'h00;
reg_space[8093] = 8'h00;
reg_space[8094] = 8'h00;
reg_space[8095] = 8'h00;
reg_space[8096] = 8'h00;
reg_space[8097] = 8'h00;
reg_space[8098] = 8'h00;
reg_space[8099] = 8'h00;
reg_space[8100; = 8'h00;
reg_space[8101] = 8'h00;
reg_space[8102] = 8'h00;
reg_space[8103] = 8'h00;
reg_space[8104] = 8'h00;
reg_space[8105] = 8'h00;
reg_space[8106] = 8'h00;
reg_space[8107] = 8'h00;
reg_space[8108] = 8'h00;
reg_space[8109] = 8'h00;
reg_space[8110] = 8'h00;
reg_space[8111] = 8'h00;
reg_space[8112] = 8'h00;
reg_space[8113] = 8'h00;
reg_space[8114] = 8'h00;
reg_space[8115] = 8'h00;
reg_space[8116] = 8'h00;
reg_space[8117] = 8'h00;
reg_space[8118] = 8'h00;
reg_space[8119] = 8'h00;
reg_space[8120] = 8'h00;
reg_space[8121] = 8'h00;
reg_space[8122] = 8'h00;
reg_space[8123] = 8'h00;
reg_space[8124] = 8'h00;
reg_space[8125] = 8'h00;
reg_space[8126] = 8'h00;
reg_space[8127] = 8'h00;
reg_space[8128] = 8'h00;
reg_space[8129] = 8'h00;
reg_space[8130] = 8'h00;
reg_space[8131] = 8'h00;
reg_space[8132] = 8'h00;
reg_space[8133] = 8'h00;
reg_space[8134] = 8'h00;
reg_space[8135] = 8'h00;
reg_space[8136] = 8'h00;
reg_space[8137] = 8'h00;
reg_space[8138] = 8'h00;
reg_space[8139] = 8'h00;
reg_space[8140] = 8'h00;
reg_space[8141] = 8'h00;
reg_space[8142] = 8'h00;
reg_space[8143] = 8'h00;
reg_space[8144] = 8'h00;
reg_space[8145] = 8'h00;
reg_space[8146] = 8'h00;
reg_space[8147] = 8'h00;
reg_space[8148] = 8'h00;
reg_space[8149] = 8'h00;
reg_space[8150] = 8'h00;
reg_space[8151] = 8'h00;
reg_space[8152] = 8'h00;
reg_space[8153] = 8'h00;
reg_space[8154] = 8'h00;
reg_space[8155] = 8'h00;
reg_space[8156] = 8'h00;
reg_space[8157] = 8'h00;
reg_space[8158] = 8'h00;
reg_space[8159] = 8'h00;
reg_space[8160] = 8'h00;
reg_space[8161] = 8'h00;
reg_space[8162] = 8'h00;
reg_space[8163] = 8'h00;
reg_space[8164] = 8'h00;
reg_space[8165] = 8'h00;
reg_space[8166] = 8'h00;
reg_space[8167] = 8'h00;
reg_space[8168] = 8'h00;
reg_space[8169] = 8'h00;
reg_space[8170] = 8'h00;
reg_space[8171] = 8'h00;
reg_space[8172] = 8'h00;
reg_space[8173] = 8'h00;
reg_space[8174] = 8'h00;
reg_space[8175] = 8'h00;
reg_space[8176] = 8'h00;
reg_space[8177] = 8'h00;
reg_space[8178] = 8'h00;
reg_space[8179] = 8'h00;
reg_space[8180] = 8'h00;
reg_space[8181] = 8'h00;
reg_space[8182] = 8'h00;
reg_space[8183] = 8'h00;
reg_space[8184] = 8'h00;
reg_space[8185] = 8'h00;
reg_space[8186] = 8'h00;
reg_space[8187] = 8'h00;
reg_space[8188] = 8'h00;
reg_space[8189] = 8'h00;
reg_space[8190] = 8'h00;
reg_space[8191] = 8'h00;
end