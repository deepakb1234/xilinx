always@(posedge ck)
begin
if(!reset || cs)
begin
maxvy_reg[512] <= 32'h00;
maxvy_reg[513] <= 32'h00;
maxvy_reg[514] <= 32'h00;
maxvy_reg[515] <= 32'h00;
maxvy_reg[516] <= 32'h00;
maxvy_reg[517] <= 32'h00;
maxvy_reg[518] <= 32'h00;
maxvy_reg[519] <= 32'h00;
maxvy_reg[520] <= 32'h00;
maxvy_reg[521] <= 32'h00;
maxvy_reg[522] <= 32'h00;
maxvy_reg[523] <= 32'h00;
maxvy_reg[524] <= 32'h00;
maxvy_reg[525] <= 32'h00;
maxvy_reg[526] <= 32'h00;
maxvy_reg[527] <= 32'h00;
maxvy_reg[528] <= 32'h00;
maxvy_reg[529] <= 32'h00;
maxvy_reg[530] <= 32'h00;
maxvy_reg[531] <= 32'h00;
maxvy_reg[532] <= 32'h00;
maxvy_reg[533] <= 32'h00;
maxvy_reg[534] <= 32'h00;
maxvy_reg[535] <= 32'h00;
maxvy_reg[536] <= 32'h00;
maxvy_reg[537] <= 32'h00;
maxvy_reg[538] <= 32'h00;
maxvy_reg[539] <= 32'h00;
maxvy_reg[540] <= 32'h00;
maxvy_reg[541] <= 32'h00;
maxvy_reg[542] <= 32'h00;
maxvy_reg[543] <= 32'h00;
maxvy_reg[544] <= 32'h00;
maxvy_reg[545] <= 32'h00;
maxvy_reg[546] <= 32'h00;
maxvy_reg[547] <= 32'h00;
maxvy_reg[548] <= 32'h00;
maxvy_reg[549] <= 32'h00;
maxvy_reg[550] <= 32'h00;
maxvy_reg[551] <= 32'h00;
maxvy_reg[552] <= 32'h00;
maxvy_reg[553] <= 32'h00;
maxvy_reg[554] <= 32'h00;
maxvy_reg[555] <= 32'h00;
maxvy_reg[556] <= 32'h00;
maxvy_reg[557] <= 32'h00;
maxvy_reg[558] <= 32'h00;
maxvy_reg[559] <= 32'h00;
maxvy_reg[560] <= 32'h00;
maxvy_reg[561] <= 32'h00;
maxvy_reg[562] <= 32'h00;
maxvy_reg[563] <= 32'h00;
maxvy_reg[564] <= 32'h00;
maxvy_reg[565] <= 32'h00;
maxvy_reg[566] <= 32'h00;
maxvy_reg[567] <= 32'h00;
maxvy_reg[568] <= 32'h00;
maxvy_reg[569] <= 32'h00;
maxvy_reg[570] <= 32'h00;
maxvy_reg[571] <= 32'h00;
maxvy_reg[572] <= 32'h00;
maxvy_reg[573] <= 32'h00;
maxvy_reg[574] <= 32'h00;
maxvy_reg[575] <= 32'h00;
maxvy_reg[576] <= 32'h00;
maxvy_reg[577] <= 32'h00;
maxvy_reg[578] <= 32'h00;
maxvy_reg[579] <= 32'h00;
maxvy_reg[580] <= 32'h00;
maxvy_reg[581] <= 32'h00;
maxvy_reg[582] <= 32'h00;
maxvy_reg[583] <= 32'h00;
maxvy_reg[584] <= 32'h00;
maxvy_reg[585] <= 32'h00;
maxvy_reg[586] <= 32'h00;
maxvy_reg[587] <= 32'h00;
maxvy_reg[588] <= 32'h00;
maxvy_reg[589] <= 32'h00;
maxvy_reg[590] <= 32'h00;
maxvy_reg[591] <= 32'h00;
maxvy_reg[592] <= 32'h00;
maxvy_reg[593] <= 32'h00;
maxvy_reg[594] <= 32'h00;
maxvy_reg[595] <= 32'h00;
maxvy_reg[596] <= 32'h00;
maxvy_reg[597] <= 32'h00;
maxvy_reg[598] <= 32'h00;
maxvy_reg[599] <= 32'h00;
maxvy_reg[600] <= 32'h00;
maxvy_reg[601] <= 32'h00;
maxvy_reg[602] <= 32'h00;
maxvy_reg[603] <= 32'h00;
maxvy_reg[604] <= 32'h00;
maxvy_reg[605] <= 32'h00;
maxvy_reg[606] <= 32'h00;
maxvy_reg[607] <= 32'h00;
maxvy_reg[608] <= 32'h00;
maxvy_reg[609] <= 32'h00;
maxvy_reg[610] <= 32'h00;
maxvy_reg[611] <= 32'h00;
maxvy_reg[612] <= 32'h00;
maxvy_reg[613] <= 32'h00;
maxvy_reg[614] <= 32'h00;
maxvy_reg[615] <= 32'h00;
maxvy_reg[616] <= 32'h00;
maxvy_reg[617] <= 32'h00;
maxvy_reg[618] <= 32'h00;
maxvy_reg[619] <= 32'h00;
maxvy_reg[620] <= 32'h00;
maxvy_reg[621] <= 32'h00;
maxvy_reg[622] <= 32'h00;
maxvy_reg[623] <= 32'h00;
maxvy_reg[624] <= 32'h00;
maxvy_reg[625] <= 32'h00;
maxvy_reg[626] <= 32'h00;
maxvy_reg[627] <= 32'h00;
maxvy_reg[628] <= 32'h00;
maxvy_reg[629] <= 32'h00;
maxvy_reg[630] <= 32'h00;
maxvy_reg[631] <= 32'h00;
maxvy_reg[632] <= 32'h00;
maxvy_reg[633] <= 32'h00;
maxvy_reg[634] <= 32'h00;
maxvy_reg[635] <= 32'h00;
maxvy_reg[636] <= 32'h00;
maxvy_reg[637] <= 32'h00;
maxvy_reg[638] <= 32'h00;
maxvy_reg[639] <= 32'h00;
maxvy_reg[640] <= 32'h00;
maxvy_reg[641] <= 32'h00;
maxvy_reg[642] <= 32'h00;
maxvy_reg[643] <= 32'h00;
maxvy_reg[644] <= 32'h00;
maxvy_reg[645] <= 32'h00;
maxvy_reg[646] <= 32'h00;
maxvy_reg[647] <= 32'h00;
maxvy_reg[648] <= 32'h00;
maxvy_reg[649] <= 32'h00;
maxvy_reg[650] <= 32'h00;
maxvy_reg[651] <= 32'h00;
maxvy_reg[652] <= 32'h00;
maxvy_reg[653] <= 32'h00;
maxvy_reg[654] <= 32'h00;
maxvy_reg[655] <= 32'h00;
maxvy_reg[656] <= 32'h00;
maxvy_reg[657] <= 32'h00;
maxvy_reg[658] <= 32'h00;
maxvy_reg[659] <= 32'h00;
maxvy_reg[660] <= 32'h00;
maxvy_reg[661] <= 32'h00;
maxvy_reg[662] <= 32'h00;
maxvy_reg[663] <= 32'h00;
maxvy_reg[664] <= 32'h00;
maxvy_reg[665] <= 32'h00;
maxvy_reg[666] <= 32'h00;
maxvy_reg[667] <= 32'h00;
maxvy_reg[668] <= 32'h00;
maxvy_reg[669] <= 32'h00;
maxvy_reg[670] <= 32'h00;
maxvy_reg[671] <= 32'h00;
maxvy_reg[672] <= 32'h00;
maxvy_reg[673] <= 32'h00;
maxvy_reg[674] <= 32'h00;
maxvy_reg[675] <= 32'h00;
maxvy_reg[676] <= 32'h00;
maxvy_reg[677] <= 32'h00;
maxvy_reg[678] <= 32'h00;
maxvy_reg[679] <= 32'h00;
maxvy_reg[680] <= 32'h00;
maxvy_reg[681] <= 32'h00;
maxvy_reg[682] <= 32'h00;
maxvy_reg[683] <= 32'h00;
maxvy_reg[684] <= 32'h00;
maxvy_reg[685] <= 32'h00;
maxvy_reg[686] <= 32'h00;
maxvy_reg[687] <= 32'h00;
maxvy_reg[688] <= 32'h00;
maxvy_reg[689] <= 32'h00;
maxvy_reg[690] <= 32'h00;
maxvy_reg[691] <= 32'h00;
maxvy_reg[692] <= 32'h00;
maxvy_reg[693] <= 32'h00;
maxvy_reg[694] <= 32'h00;
maxvy_reg[695] <= 32'h00;
maxvy_reg[696] <= 32'h00;
maxvy_reg[697] <= 32'h00;
maxvy_reg[698] <= 32'h00;
maxvy_reg[699] <= 32'h00;
maxvy_reg[700] <= 32'h00;
maxvy_reg[701] <= 32'h00;
maxvy_reg[702] <= 32'h00;
maxvy_reg[703] <= 32'h00;
maxvy_reg[704] <= 32'h00;
maxvy_reg[705] <= 32'h00;
maxvy_reg[706] <= 32'h00;
maxvy_reg[707] <= 32'h00;
maxvy_reg[708] <= 32'h00;
maxvy_reg[709] <= 32'h00;
maxvy_reg[710] <= 32'h00;
maxvy_reg[711] <= 32'h00;
maxvy_reg[712] <= 32'h00;
maxvy_reg[713] <= 32'h00;
maxvy_reg[714] <= 32'h00;
maxvy_reg[715] <= 32'h00;
maxvy_reg[716] <= 32'h00;
maxvy_reg[717] <= 32'h00;
maxvy_reg[718] <= 32'h00;
maxvy_reg[719] <= 32'h00;
maxvy_reg[720] <= 32'h00;
maxvy_reg[721] <= 32'h00;
maxvy_reg[722] <= 32'h00;
maxvy_reg[723] <= 32'h00;
maxvy_reg[724] <= 32'h00;
maxvy_reg[725] <= 32'h00;
maxvy_reg[726] <= 32'h00;
maxvy_reg[727] <= 32'h00;
maxvy_reg[728] <= 32'h00;
maxvy_reg[729] <= 32'h00;
maxvy_reg[730] <= 32'h00;
maxvy_reg[731] <= 32'h00;
maxvy_reg[732] <= 32'h00;
maxvy_reg[733] <= 32'h00;
maxvy_reg[734] <= 32'h00;
maxvy_reg[735] <= 32'h00;
maxvy_reg[736] <= 32'h00;
maxvy_reg[737] <= 32'h00;
maxvy_reg[738] <= 32'h00;
maxvy_reg[739] <= 32'h00;
maxvy_reg[740] <= 32'h00;
maxvy_reg[741] <= 32'h00;
maxvy_reg[742] <= 32'h00;
maxvy_reg[743] <= 32'h00;
maxvy_reg[744] <= 32'h00;
maxvy_reg[745] <= 32'h00;
maxvy_reg[746] <= 32'h00;
maxvy_reg[747] <= 32'h00;
maxvy_reg[748] <= 32'h00;
maxvy_reg[749] <= 32'h00;
maxvy_reg[750] <= 32'h00;
maxvy_reg[751] <= 32'h00;
maxvy_reg[752] <= 32'h00;
maxvy_reg[753] <= 32'h00;
maxvy_reg[754] <= 32'h00;
maxvy_reg[755] <= 32'h00;
maxvy_reg[756] <= 32'h00;
maxvy_reg[757] <= 32'h00;
maxvy_reg[758] <= 32'h00;
maxvy_reg[759] <= 32'h00;
maxvy_reg[760] <= 32'h00;
maxvy_reg[761] <= 32'h00;
maxvy_reg[762] <= 32'h00;
maxvy_reg[763] <= 32'h00;
maxvy_reg[764] <= 32'h00;
maxvy_reg[765] <= 32'h00;
maxvy_reg[766] <= 32'h00;
maxvy_reg[767] <= 32'h00;
end
else if(sdr_en && data_cnt>0 && ns==READ_DATA && command_code==32'h7F)
begin
maxvy_reg[comm_addr_reg[9:0]+{2'd0,sdr_count}][(bit_count[2:0])] <= rd_data[0];
//maxvy_reg[comm_addr_reg[31:0]][((addr_cnt-1)*8)+bit_count[2:0]] <= rd_data[0];
end
else
begin
maxvy_reg[512] <= 32'h00;
maxvy_reg[513] <= 32'h00;
maxvy_reg[514] <= 32'h00;
maxvy_reg[515] <= 32'h00;
maxvy_reg[516] <= 32'h00;
maxvy_reg[517] <= 32'h00;
maxvy_reg[518] <= 32'h00;
maxvy_reg[519] <= 32'h00;
maxvy_reg[520] <= 32'h00;
maxvy_reg[521] <= 32'h00;
maxvy_reg[522] <= 32'h00;
maxvy_reg[523] <= 32'h00;
maxvy_reg[524] <= 32'h00;
maxvy_reg[525] <= 32'h00;
maxvy_reg[526] <= 32'h00;
maxvy_reg[527] <= 32'h00;
maxvy_reg[528] <= 32'h00;
maxvy_reg[529] <= 32'h00;
maxvy_reg[530] <= 32'h00;
maxvy_reg[531] <= 32'h00;
maxvy_reg[532] <= 32'h00;
maxvy_reg[533] <= 32'h00;
maxvy_reg[534] <= 32'h00;
maxvy_reg[535] <= 32'h00;
maxvy_reg[536] <= 32'h00;
maxvy_reg[537] <= 32'h00;
maxvy_reg[538] <= 32'h00;
maxvy_reg[539] <= 32'h00;
maxvy_reg[540] <= 32'h00;
maxvy_reg[541] <= 32'h00;
maxvy_reg[542] <= 32'h00;
maxvy_reg[543] <= 32'h00;
maxvy_reg[544] <= 32'h00;
maxvy_reg[545] <= 32'h00;
maxvy_reg[546] <= 32'h00;
maxvy_reg[547] <= 32'h00;
maxvy_reg[548] <= 32'h00;
maxvy_reg[549] <= 32'h00;
maxvy_reg[550] <= 32'h00;
maxvy_reg[551] <= 32'h00;
maxvy_reg[552] <= 32'h00;
maxvy_reg[553] <= 32'h00;
maxvy_reg[554] <= 32'h00;
maxvy_reg[555] <= 32'h00;
maxvy_reg[556] <= 32'h00;
maxvy_reg[557] <= 32'h00;
maxvy_reg[558] <= 32'h00;
maxvy_reg[559] <= 32'h00;
maxvy_reg[560] <= 32'h00;
maxvy_reg[561] <= 32'h00;
maxvy_reg[562] <= 32'h00;
maxvy_reg[563] <= 32'h00;
maxvy_reg[564] <= 32'h00;
maxvy_reg[565] <= 32'h00;
maxvy_reg[566] <= 32'h00;
maxvy_reg[567] <= 32'h00;
maxvy_reg[568] <= 32'h00;
maxvy_reg[569] <= 32'h00;
maxvy_reg[570] <= 32'h00;
maxvy_reg[571] <= 32'h00;
maxvy_reg[572] <= 32'h00;
maxvy_reg[573] <= 32'h00;
maxvy_reg[574] <= 32'h00;
maxvy_reg[575] <= 32'h00;
maxvy_reg[576] <= 32'h00;
maxvy_reg[577] <= 32'h00;
maxvy_reg[578] <= 32'h00;
maxvy_reg[579] <= 32'h00;
maxvy_reg[580] <= 32'h00;
maxvy_reg[581] <= 32'h00;
maxvy_reg[582] <= 32'h00;
maxvy_reg[583] <= 32'h00;
maxvy_reg[584] <= 32'h00;
maxvy_reg[585] <= 32'h00;
maxvy_reg[586] <= 32'h00;
maxvy_reg[587] <= 32'h00;
maxvy_reg[588] <= 32'h00;
maxvy_reg[589] <= 32'h00;
maxvy_reg[590] <= 32'h00;
maxvy_reg[591] <= 32'h00;
maxvy_reg[592] <= 32'h00;
maxvy_reg[593] <= 32'h00;
maxvy_reg[594] <= 32'h00;
maxvy_reg[595] <= 32'h00;
maxvy_reg[596] <= 32'h00;
maxvy_reg[597] <= 32'h00;
maxvy_reg[598] <= 32'h00;
maxvy_reg[599] <= 32'h00;
maxvy_reg[600] <= 32'h00;
maxvy_reg[601] <= 32'h00;
maxvy_reg[602] <= 32'h00;
maxvy_reg[603] <= 32'h00;
maxvy_reg[604] <= 32'h00;
maxvy_reg[605] <= 32'h00;
maxvy_reg[606] <= 32'h00;
maxvy_reg[607] <= 32'h00;
maxvy_reg[608] <= 32'h00;
maxvy_reg[609] <= 32'h00;
maxvy_reg[610] <= 32'h00;
maxvy_reg[611] <= 32'h00;
maxvy_reg[612] <= 32'h00;
maxvy_reg[613] <= 32'h00;
maxvy_reg[614] <= 32'h00;
maxvy_reg[615] <= 32'h00;
maxvy_reg[616] <= 32'h00;
maxvy_reg[617] <= 32'h00;
maxvy_reg[618] <= 32'h00;
maxvy_reg[619] <= 32'h00;
maxvy_reg[620] <= 32'h00;
maxvy_reg[621] <= 32'h00;
maxvy_reg[622] <= 32'h00;
maxvy_reg[623] <= 32'h00;
maxvy_reg[624] <= 32'h00;
maxvy_reg[625] <= 32'h00;
maxvy_reg[626] <= 32'h00;
maxvy_reg[627] <= 32'h00;
maxvy_reg[628] <= 32'h00;
maxvy_reg[629] <= 32'h00;
maxvy_reg[630] <= 32'h00;
maxvy_reg[631] <= 32'h00;
maxvy_reg[632] <= 32'h00;
maxvy_reg[633] <= 32'h00;
maxvy_reg[634] <= 32'h00;
maxvy_reg[635] <= 32'h00;
maxvy_reg[636] <= 32'h00;
maxvy_reg[637] <= 32'h00;
maxvy_reg[638] <= 32'h00;
maxvy_reg[639] <= 32'h00;
maxvy_reg[640] <= 32'h00;
maxvy_reg[641] <= 32'h00;
maxvy_reg[642] <= 32'h00;
maxvy_reg[643] <= 32'h00;
maxvy_reg[644] <= 32'h00;
maxvy_reg[645] <= 32'h00;
maxvy_reg[646] <= 32'h00;
maxvy_reg[647] <= 32'h00;
maxvy_reg[648] <= 32'h00;
maxvy_reg[649] <= 32'h00;
maxvy_reg[650] <= 32'h00;
maxvy_reg[651] <= 32'h00;
maxvy_reg[652] <= 32'h00;
maxvy_reg[653] <= 32'h00;
maxvy_reg[654] <= 32'h00;
maxvy_reg[655] <= 32'h00;
maxvy_reg[656] <= 32'h00;
maxvy_reg[657] <= 32'h00;
maxvy_reg[658] <= 32'h00;
maxvy_reg[659] <= 32'h00;
maxvy_reg[660] <= 32'h00;
maxvy_reg[661] <= 32'h00;
maxvy_reg[662] <= 32'h00;
maxvy_reg[663] <= 32'h00;
maxvy_reg[664] <= 32'h00;
maxvy_reg[665] <= 32'h00;
maxvy_reg[666] <= 32'h00;
maxvy_reg[667] <= 32'h00;
maxvy_reg[668] <= 32'h00;
maxvy_reg[669] <= 32'h00;
maxvy_reg[670] <= 32'h00;
maxvy_reg[671] <= 32'h00;
maxvy_reg[672] <= 32'h00;
maxvy_reg[673] <= 32'h00;
maxvy_reg[674] <= 32'h00;
maxvy_reg[675] <= 32'h00;
maxvy_reg[676] <= 32'h00;
maxvy_reg[677] <= 32'h00;
maxvy_reg[678] <= 32'h00;
maxvy_reg[679] <= 32'h00;
maxvy_reg[680] <= 32'h00;
maxvy_reg[681] <= 32'h00;
maxvy_reg[682] <= 32'h00;
maxvy_reg[683] <= 32'h00;
maxvy_reg[684] <= 32'h00;
maxvy_reg[685] <= 32'h00;
maxvy_reg[686] <= 32'h00;
maxvy_reg[687] <= 32'h00;
maxvy_reg[688] <= 32'h00;
maxvy_reg[689] <= 32'h00;
maxvy_reg[690] <= 32'h00;
maxvy_reg[691] <= 32'h00;
maxvy_reg[692] <= 32'h00;
maxvy_reg[693] <= 32'h00;
maxvy_reg[694] <= 32'h00;
maxvy_reg[695] <= 32'h00;
maxvy_reg[696] <= 32'h00;
maxvy_reg[697] <= 32'h00;
maxvy_reg[698] <= 32'h00;
maxvy_reg[699] <= 32'h00;
maxvy_reg[700] <= 32'h00;
maxvy_reg[701] <= 32'h00;
maxvy_reg[702] <= 32'h00;
maxvy_reg[703] <= 32'h00;
maxvy_reg[704] <= 32'h00;
maxvy_reg[705] <= 32'h00;
maxvy_reg[706] <= 32'h00;
maxvy_reg[707] <= 32'h00;
maxvy_reg[708] <= 32'h00;
maxvy_reg[709] <= 32'h00;
maxvy_reg[710] <= 32'h00;
maxvy_reg[711] <= 32'h00;
maxvy_reg[712] <= 32'h00;
maxvy_reg[713] <= 32'h00;
maxvy_reg[714] <= 32'h00;
maxvy_reg[715] <= 32'h00;
maxvy_reg[716] <= 32'h00;
maxvy_reg[717] <= 32'h00;
maxvy_reg[718] <= 32'h00;
maxvy_reg[719] <= 32'h00;
maxvy_reg[720] <= 32'h00;
maxvy_reg[721] <= 32'h00;
maxvy_reg[722] <= 32'h00;
maxvy_reg[723] <= 32'h00;
maxvy_reg[724] <= 32'h00;
maxvy_reg[725] <= 32'h00;
maxvy_reg[726] <= 32'h00;
maxvy_reg[727] <= 32'h00;
maxvy_reg[728] <= 32'h00;
maxvy_reg[729] <= 32'h00;
maxvy_reg[730] <= 32'h00;
maxvy_reg[731] <= 32'h00;
maxvy_reg[732] <= 32'h00;
maxvy_reg[733] <= 32'h00;
maxvy_reg[734] <= 32'h00;
maxvy_reg[735] <= 32'h00;
maxvy_reg[736] <= 32'h00;
maxvy_reg[737] <= 32'h00;
maxvy_reg[738] <= 32'h00;
maxvy_reg[739] <= 32'h00;
maxvy_reg[740] <= 32'h00;
maxvy_reg[741] <= 32'h00;
maxvy_reg[742] <= 32'h00;
maxvy_reg[743] <= 32'h00;
maxvy_reg[744] <= 32'h00;
maxvy_reg[745] <= 32'h00;
maxvy_reg[746] <= 32'h00;
maxvy_reg[747] <= 32'h00;
maxvy_reg[748] <= 32'h00;
maxvy_reg[749] <= 32'h00;
maxvy_reg[750] <= 32'h00;
maxvy_reg[751] <= 32'h00;
maxvy_reg[752] <= 32'h00;
maxvy_reg[753] <= 32'h00;
maxvy_reg[754] <= 32'h00;
maxvy_reg[755] <= 32'h00;
maxvy_reg[756] <= 32'h00;
maxvy_reg[757] <= 32'h00;
maxvy_reg[758] <= 32'h00;
maxvy_reg[759] <= 32'h00;
maxvy_reg[760] <= 32'h00;
maxvy_reg[761] <= 32'h00;
maxvy_reg[762] <= 32'h00;
maxvy_reg[763] <= 32'h00;
maxvy_reg[764] <= 32'h00;
maxvy_reg[765] <= 32'h00;
maxvy_reg[766] <= 32'h00;
maxvy_reg[767] <= 32'h00;
end
end