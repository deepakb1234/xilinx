always@(reset)
begin
 
	sfdp_hdr_reg[0]=8'h53;
	sfdp_hdr_reg[1]=8'h46;
	sfdp_hdr_reg[2]=8'h44;
	sfdp_hdr_reg[3]=8'h50;

	sfdp_hdr_reg[4]=8'h00;
	sfdp_hdr_reg[5]=8'h01;
	sfdp_hdr_reg[6]=8'h00;
	sfdp_hdr_reg[7]=8'hFA;

	sfdp_hdr_reg[8]=8'h06;
	sfdp_hdr_reg[9]=8'h00;
	sfdp_hdr_reg[10]=8'h01;
	sfdp_hdr_reg[11]=8'h08;

	sfdp_hdr_reg[12]=8'h30;
	sfdp_hdr_reg[13]=8'h00;
	sfdp_hdr_reg[14]=8'h00;
	sfdp_hdr_reg[15]=8'hFF;

	sfdp_hdr_reg[16]=8'h06;
	sfdp_hdr_reg[17]=8'h00;
	sfdp_hdr_reg[18]=8'h01;
	sfdp_hdr_reg[19]=8'h09;

	sfdp_hdr_reg[20]=8'h60;
	sfdp_hdr_reg[21]=8'h00;
	sfdp_hdr_reg[22]=8'h00;
	sfdp_hdr_reg[23]=8'hFF;

//*******SFDP PARAMETER REGISTER*********//
	sfdp_hdr_reg[24]=8'hE0;
	sfdp_hdr_reg[25]=8'hFF;
	sfdp_hdr_reg[26]=8'hFF;
	sfdp_hdr_reg[27]=8'hFF;

	sfdp_hdr_reg[28]=8'h10;
	sfdp_hdr_reg[29]=8'h02;
	sfdp_hdr_reg[30]=8'h00;
	sfdp_hdr_reg[31]=8'h00;

	sfdp_hdr_reg[32]=8'h00;
	sfdp_hdr_reg[33]=8'h00;
	sfdp_hdr_reg[34]=8'h00;
	sfdp_hdr_reg[35]=8'h00;
sfdp_hdr_reg[36] = 8'h00;
sfdp_hdr_reg[37] = 8'h00;
sfdp_hdr_reg[38] = 8'h00;
sfdp_hdr_reg[39] = 8'h00;
sfdp_hdr_reg[40] = 8'h00;
sfdp_hdr_reg[41] = 8'h00;
sfdp_hdr_reg[42] = 8'h00;
sfdp_hdr_reg[43] = 8'h00;
sfdp_hdr_reg[44] = 8'h00;
sfdp_hdr_reg[45] = 8'h00;
sfdp_hdr_reg[46] = 8'h00;
sfdp_hdr_reg[47] = 8'h00;
sfdp_hdr_reg[48] = 8'h00;
sfdp_hdr_reg[49] = 8'h00;
sfdp_hdr_reg[50] = 8'h00;
sfdp_hdr_reg[51] = 8'h00;
sfdp_hdr_reg[52] = 8'h00;
sfdp_hdr_reg[53] = 8'h00;
sfdp_hdr_reg[54] = 8'h00;
sfdp_hdr_reg[55] = 8'h00;
sfdp_hdr_reg[56] = 8'h00;
sfdp_hdr_reg[57] = 8'h00;
sfdp_hdr_reg[58] = 8'h00;
sfdp_hdr_reg[59] = 8'h00;
sfdp_hdr_reg[60] = 8'h00;
sfdp_hdr_reg[61] = 8'h00;
sfdp_hdr_reg[62] = 8'h00;
sfdp_hdr_reg[63] = 8'h00;
sfdp_hdr_reg[64] = 8'h00;
sfdp_hdr_reg[65] = 8'h00;
sfdp_hdr_reg[66] = 8'h00;
sfdp_hdr_reg[67] = 8'h00;
sfdp_hdr_reg[68] = 8'h00;
sfdp_hdr_reg[69] = 8'h00;
sfdp_hdr_reg[70] = 8'h00;
sfdp_hdr_reg[71] = 8'h00;
sfdp_hdr_reg[72] = 8'h00;
sfdp_hdr_reg[73] = 8'h00;
sfdp_hdr_reg[74] = 8'h00;
sfdp_hdr_reg[75] = 8'h00;
sfdp_hdr_reg[76] = 8'h00;
sfdp_hdr_reg[77] = 8'h00;
sfdp_hdr_reg[78] = 8'h00;
sfdp_hdr_reg[79] = 8'h00;
sfdp_hdr_reg[80] = 8'h00;
sfdp_hdr_reg[81] = 8'h00;
sfdp_hdr_reg[82] = 8'h00;
sfdp_hdr_reg[83] = 8'h00;
sfdp_hdr_reg[84] = 8'h00;
sfdp_hdr_reg[85] = 8'h00;
sfdp_hdr_reg[86] = 8'h00;
sfdp_hdr_reg[87] = 8'h00;
sfdp_hdr_reg[88] = 8'h00;
sfdp_hdr_reg[89] = 8'h00;
sfdp_hdr_reg[90] = 8'h00;
sfdp_hdr_reg[91] = 8'h00;
sfdp_hdr_reg[92] = 8'h00;
sfdp_hdr_reg[93] = 8'h00;
sfdp_hdr_reg[94] = 8'h00;
sfdp_hdr_reg[95] = 8'h00;
sfdp_hdr_reg[96] = 8'h00;
sfdp_hdr_reg[97] = 8'h00;
sfdp_hdr_reg[98] = 8'h00;
sfdp_hdr_reg[99] = 8'h00;
sfdp_hdr_reg[100] = 8'h00;
sfdp_hdr_reg[101] = 8'h00;
sfdp_hdr_reg[102] = 8'h00;
sfdp_hdr_reg[103] = 8'h00;
sfdp_hdr_reg[104] = 8'h00;
sfdp_hdr_reg[105] = 8'h00;
sfdp_hdr_reg[106] = 8'h00;
sfdp_hdr_reg[107] = 8'h00;
sfdp_hdr_reg[108] = 8'h00;
sfdp_hdr_reg[109] = 8'h00;
sfdp_hdr_reg[110] = 8'h00;
sfdp_hdr_reg[111] = 8'h00;
sfdp_hdr_reg[112] = 8'h00;
sfdp_hdr_reg[113] = 8'h00;
sfdp_hdr_reg[114] = 8'h00;
sfdp_hdr_reg[115] = 8'h00;
sfdp_hdr_reg[116] = 8'h00;
sfdp_hdr_reg[117] = 8'h00;
sfdp_hdr_reg[118] = 8'h00;
sfdp_hdr_reg[119] = 8'h00;
sfdp_hdr_reg[120] = 8'h00;
sfdp_hdr_reg[121] = 8'h00;
sfdp_hdr_reg[122] = 8'h00;
sfdp_hdr_reg[123] = 8'h00;
sfdp_hdr_reg[124] = 8'h00;
sfdp_hdr_reg[125] = 8'h00;
sfdp_hdr_reg[126] = 8'h00;
sfdp_hdr_reg[127] = 8'h00;
sfdp_hdr_reg[128] = 8'h00;
sfdp_hdr_reg[129] = 8'h00;
sfdp_hdr_reg[130] = 8'h00;
sfdp_hdr_reg[131] = 8'h00;
sfdp_hdr_reg[132] = 8'h00;
sfdp_hdr_reg[133] = 8'h00;
sfdp_hdr_reg[134] = 8'h00;
sfdp_hdr_reg[135] = 8'h00;
sfdp_hdr_reg[136] = 8'h00;
sfdp_hdr_reg[137] = 8'h00;
sfdp_hdr_reg[138] = 8'h00;
sfdp_hdr_reg[139] = 8'h00;
sfdp_hdr_reg[140] = 8'h00;
sfdp_hdr_reg[141] = 8'h00;
sfdp_hdr_reg[142] = 8'h00;
sfdp_hdr_reg[143] = 8'h00;
sfdp_hdr_reg[144] = 8'h00;
sfdp_hdr_reg[145] = 8'h00;
sfdp_hdr_reg[146] = 8'h00;
sfdp_hdr_reg[147] = 8'h00;
sfdp_hdr_reg[148] = 8'h00;
sfdp_hdr_reg[149] = 8'h00;
sfdp_hdr_reg[150] = 8'h00;
sfdp_hdr_reg[151] = 8'h00;
sfdp_hdr_reg[152] = 8'h00;
sfdp_hdr_reg[153] = 8'h00;
sfdp_hdr_reg[154] = 8'h00;
sfdp_hdr_reg[155] = 8'h00;
sfdp_hdr_reg[156] = 8'h00;
sfdp_hdr_reg[157] = 8'h00;
sfdp_hdr_reg[158] = 8'h00;
sfdp_hdr_reg[159] = 8'h00;
sfdp_hdr_reg[160] = 8'h00;
sfdp_hdr_reg[161] = 8'h00;
sfdp_hdr_reg[162] = 8'h00;
sfdp_hdr_reg[163] = 8'h00;
sfdp_hdr_reg[164] = 8'h00;
sfdp_hdr_reg[165] = 8'h00;
sfdp_hdr_reg[166] = 8'h00;
sfdp_hdr_reg[167] = 8'h00;
sfdp_hdr_reg[168] = 8'h00;
sfdp_hdr_reg[169] = 8'h00;
sfdp_hdr_reg[170] = 8'h00;
sfdp_hdr_reg[171] = 8'h00;
sfdp_hdr_reg[172] = 8'h00;
sfdp_hdr_reg[173] = 8'h00;
sfdp_hdr_reg[174] = 8'h00;
sfdp_hdr_reg[175] = 8'h00;
sfdp_hdr_reg[176] = 8'h00;
sfdp_hdr_reg[177] = 8'h00;
sfdp_hdr_reg[178] = 8'h00;
sfdp_hdr_reg[179] = 8'h00;
sfdp_hdr_reg[180] = 8'h00;
sfdp_hdr_reg[181] = 8'h00;
sfdp_hdr_reg[182] = 8'h00;
sfdp_hdr_reg[183] = 8'h00;
sfdp_hdr_reg[184] = 8'h00;
sfdp_hdr_reg[185] = 8'h00;
sfdp_hdr_reg[186] = 8'h00;
sfdp_hdr_reg[187] = 8'h00;
sfdp_hdr_reg[188] = 8'h00;
sfdp_hdr_reg[189] = 8'h00;
sfdp_hdr_reg[190] = 8'h00;
sfdp_hdr_reg[191] = 8'h00;
sfdp_hdr_reg[192] = 8'h00;
sfdp_hdr_reg[193] = 8'h00;
sfdp_hdr_reg[194] = 8'h00;
sfdp_hdr_reg[195] = 8'h00;
sfdp_hdr_reg[196] = 8'h00;
sfdp_hdr_reg[197] = 8'h00;
sfdp_hdr_reg[198] = 8'h00;
sfdp_hdr_reg[199] = 8'h00;
sfdp_hdr_reg[200] = 8'h00;
sfdp_hdr_reg[201] = 8'h00;
sfdp_hdr_reg[202] = 8'h00;
sfdp_hdr_reg[203] = 8'h00;
sfdp_hdr_reg[204] = 8'h00;
sfdp_hdr_reg[205] = 8'h00;
sfdp_hdr_reg[206] = 8'h00;
sfdp_hdr_reg[207] = 8'h00;
sfdp_hdr_reg[208] = 8'h00;
sfdp_hdr_reg[209] = 8'h00;
sfdp_hdr_reg[210] = 8'h00;
sfdp_hdr_reg[211] = 8'h00;
sfdp_hdr_reg[212] = 8'h00;
sfdp_hdr_reg[213] = 8'h00;
sfdp_hdr_reg[214] = 8'h00;
sfdp_hdr_reg[215] = 8'h00;
sfdp_hdr_reg[216] = 8'h00;
sfdp_hdr_reg[217] = 8'h00;
sfdp_hdr_reg[218] = 8'h00;
sfdp_hdr_reg[219] = 8'h00;
sfdp_hdr_reg[220] = 8'h00;
sfdp_hdr_reg[221] = 8'h00;
sfdp_hdr_reg[222] = 8'h00;
sfdp_hdr_reg[223] = 8'h00;
sfdp_hdr_reg[224] = 8'h00;
sfdp_hdr_reg[225] = 8'h00;
sfdp_hdr_reg[226] = 8'h00;
sfdp_hdr_reg[227] = 8'h00;
sfdp_hdr_reg[228] = 8'h00;
sfdp_hdr_reg[229] = 8'h00;
sfdp_hdr_reg[230] = 8'h00;
sfdp_hdr_reg[231] = 8'h00;
sfdp_hdr_reg[232] = 8'h00;
sfdp_hdr_reg[233] = 8'h00;
sfdp_hdr_reg[234] = 8'h00;
sfdp_hdr_reg[235] = 8'h00;
sfdp_hdr_reg[236] = 8'h00;
sfdp_hdr_reg[237] = 8'h00;
sfdp_hdr_reg[238] = 8'h00;
sfdp_hdr_reg[239] = 8'h00;
sfdp_hdr_reg[240] = 8'h00;
sfdp_hdr_reg[241] = 8'h00;
sfdp_hdr_reg[242] = 8'h00;
sfdp_hdr_reg[243] = 8'h00;
sfdp_hdr_reg[244] = 8'h00;
sfdp_hdr_reg[245] = 8'h00;
sfdp_hdr_reg[246] = 8'h00;
sfdp_hdr_reg[247] = 8'h00;
sfdp_hdr_reg[248] = 8'h00;
sfdp_hdr_reg[249] = 8'h00;
sfdp_hdr_reg[250] = 8'h00;
sfdp_hdr_reg[251] = 8'h00;
sfdp_hdr_reg[252] = 8'h00;
sfdp_hdr_reg[253] = 8'h00;
sfdp_hdr_reg[254] = 8'h00;
sfdp_hdr_reg[255] = 8'h00;
end
