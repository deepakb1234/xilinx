always@(reset)
begin
sccr_reg[256] = 8'h53;
	sccr_reg[257] = 8'h46;
	sccr_reg[258] = 8'h44;
	sccr_reg[259] = 8'h50;

	sccr_reg[260] = 8'h00;
	sccr_reg[261] = 8'h01;
	sccr_reg[262] = 8'h00;
	sccr_reg[263] = 8'hFA;

	sccr_reg[264] = 8'h09;
	sccr_reg[265] = 8'h00;
	sccr_reg[266] = 8'h01;
	sccr_reg[267] = 8'h08;

	sccr_reg[268] = 8'h30;
	sccr_reg[269] = 8'h00;
	sccr_reg[270] = 8'h00;
	sccr_reg[271] = 8'hFF;

	sccr_reg[272] = 8'hab;
	sccr_reg[273] = 8'hab;
	sccr_reg[274] = 8'hab;
	sccr_reg[275] = 8'hab;

	sccr_reg[276] = 8'hab;
	sccr_reg[277] = 8'hab;
	sccr_reg[278] = 8'hab;
	sccr_reg[279] = 8'hab;

	sccr_reg[280] = 8'hc2;
	sccr_reg[281] = 8'h12;
	sccr_reg[282] = 8'h98;
	sccr_reg[283] = 8'h00;

	sccr_reg[284] = 8'hb4;
	sccr_reg[285] = 8'h10;
	sccr_reg[286] = 8'h00;
	sccr_reg[287] = 8'h00;

	sccr_reg[288] = 8'hb4;
	sccr_reg[289] = 8'h10;
	sccr_reg[290] = 8'h00;
	sccr_reg[291] = 8'h00;

	sccr_reg[292] = 8'ha2;
	sccr_reg[293] = 8'h10;
	sccr_reg[294] = 8'h00;
	sccr_reg[295] = 8'h00;

	sccr_reg[296] = 8'ha2;
	sccr_reg[297] = 8'h10;
	sccr_reg[298] = 8'h00;
	sccr_reg[299] = 8'h00;

	sccr_reg[300] = 8'h92;
	sccr_reg[301] = 8'h49;
	sccr_reg[302] = 8'h24;
	sccr_reg[303] = 8'h90;

	sccr_reg[304] = 8'h92;
	sccr_reg[305] = 8'h49;
	sccr_reg[306] = 8'h24;
	sccr_reg[307] = 8'h90;

	sccr_reg[308] = 8'h92;
	sccr_reg[309] = 8'h49;
	sccr_reg[310] = 8'h24;
	sccr_reg[311] = 8'h90;

	sccr_reg[312] = 8'h68;
	sccr_reg[313] = 8'h20;
	sccr_reg[314] = 8'h00;
	sccr_reg[315] = 8'h00;

	sccr_reg[316] = 8'h68;
	sccr_reg[317] = 8'h20;
	sccr_reg[318] = 8'h00;
	sccr_reg[319] = 8'h00;
	
	
sccr_reg[320] = 8'h00;
sccr_reg[321] = 8'h00;
sccr_reg[322] = 8'h00;
sccr_reg[323] = 8'h00;
sccr_reg[324] = 8'h00;
sccr_reg[325] = 8'h00;
sccr_reg[326] = 8'h00;
sccr_reg[327] = 8'h00;
sccr_reg[328] = 8'h00;
sccr_reg[329] = 8'h00;
sccr_reg[330] = 8'h00;
sccr_reg[331] = 8'h00;
sccr_reg[332] = 8'h00;
sccr_reg[333] = 8'h00;
sccr_reg[334] = 8'h00;
sccr_reg[335] = 8'h00;
sccr_reg[336] = 8'h00;
sccr_reg[337] = 8'h00;
sccr_reg[338] = 8'h00;
sccr_reg[339] = 8'h00;
sccr_reg[340] = 8'h00;
sccr_reg[341] = 8'h00;
sccr_reg[342] = 8'h00;
sccr_reg[343] = 8'h00;
sccr_reg[344] = 8'h00;
sccr_reg[345] = 8'h00;
sccr_reg[346] = 8'h00;
sccr_reg[347] = 8'h00;
sccr_reg[348] = 8'h00;
sccr_reg[349] = 8'h00;

sccr_reg[350] = 8'h00;
sccr_reg[351] = 8'h00;
sccr_reg[352] = 8'h00;
sccr_reg[353] = 8'h00;
sccr_reg[354] = 8'h00;
sccr_reg[355] = 8'h00;
sccr_reg[356] = 8'h00;
sccr_reg[357] = 8'h00;
sccr_reg[358] = 8'h00;
sccr_reg[359] = 8'h00;

sccr_reg[360] = 8'h00;
sccr_reg[361] = 8'h00;
sccr_reg[362] = 8'h00;
sccr_reg[363] = 8'h00;
sccr_reg[364] = 8'h00;
sccr_reg[365] = 8'h00;
sccr_reg[366] = 8'h00;
sccr_reg[367] = 8'h00;
sccr_reg[368] = 8'h00;
sccr_reg[369] = 8'h00;
sccr_reg[370] = 8'h00;
sccr_reg[371] = 8'h00;
sccr_reg[372] = 8'h00;
sccr_reg[373] = 8'h00;
sccr_reg[374] = 8'h00;
sccr_reg[375] = 8'h00;
sccr_reg[376] = 8'h00;
sccr_reg[377] = 8'h00;
sccr_reg[378] = 8'h00;
sccr_reg[379] = 8'h00;
sccr_reg[380] = 8'h00;
sccr_reg[381] = 8'h00;
sccr_reg[382] = 8'h00;
sccr_reg[383] = 8'h00;
sccr_reg[384] = 8'h00;
sccr_reg[385] = 8'h00;
sccr_reg[386] = 8'h00;
sccr_reg[387] = 8'h00;
sccr_reg[388] = 8'h00;
sccr_reg[389] = 8'h00;
sccr_reg[390] = 8'h00;
sccr_reg[391] = 8'h00;
sccr_reg[392] = 8'h00;
sccr_reg[393] = 8'h00;
sccr_reg[394] = 8'h00;
sccr_reg[395] = 8'h00;
sccr_reg[396] = 8'h00;
sccr_reg[397] = 8'h00;
sccr_reg[398] = 8'h00;
sccr_reg[399] = 8'h00;
sccr_reg[400] = 8'h00;
sccr_reg[401] = 8'h00;
sccr_reg[402] = 8'h00;
sccr_reg[403] = 8'h00;
sccr_reg[404] = 8'h00;
sccr_reg[405] = 8'h00;
sccr_reg[406] = 8'h00;
sccr_reg[407] = 8'h00;
sccr_reg[408] = 8'h00;
sccr_reg[409] = 8'h00;
sccr_reg[410] = 8'h00;
sccr_reg[411] = 8'h00;
sccr_reg[412] = 8'h00;
sccr_reg[413] = 8'h00;
sccr_reg[414] = 8'h00;
sccr_reg[415] = 8'h00;
sccr_reg[416] = 8'h00;
sccr_reg[417] = 8'h00;
sccr_reg[418] = 8'h00;
sccr_reg[419] = 8'h00;
sccr_reg[420] = 8'h00;
sccr_reg[421] = 8'h00;
sccr_reg[422] = 8'h00;
sccr_reg[423] = 8'h00;
sccr_reg[424] = 8'h00;
sccr_reg[425] = 8'h00;
sccr_reg[426] = 8'h00;
sccr_reg[427] = 8'h00;
sccr_reg[428] = 8'h00;
sccr_reg[429] = 8'h00;
sccr_reg[430] = 8'h00;
sccr_reg[431] = 8'h00;
sccr_reg[432] = 8'h00;
sccr_reg[433] = 8'h00;
sccr_reg[434] = 8'h00;
sccr_reg[435] = 8'h00;
sccr_reg[436] = 8'h00;
sccr_reg[437] = 8'h00;
sccr_reg[438] = 8'h00;
sccr_reg[439] = 8'h00;
sccr_reg[440] = 8'h00;
sccr_reg[441] = 8'h00;
sccr_reg[442] = 8'h00;
sccr_reg[443] = 8'h00;
sccr_reg[444] = 8'h00;
sccr_reg[445] = 8'h00;
sccr_reg[446] = 8'h00;
sccr_reg[447] = 8'h00;
sccr_reg[448] = 8'h00;
sccr_reg[449] = 8'h00;
sccr_reg[450] = 8'h00;
sccr_reg[451] = 8'h00;
sccr_reg[452] = 8'h00;
sccr_reg[453] = 8'h00;
sccr_reg[454] = 8'h00;
sccr_reg[455] = 8'h00;
sccr_reg[456] = 8'h00;
sccr_reg[457] = 8'h00;
sccr_reg[458] = 8'h00;
sccr_reg[459] = 8'h00;
sccr_reg[460] = 8'h00;
sccr_reg[461] = 8'h00;
sccr_reg[462] = 8'h00;
sccr_reg[463] = 8'h00;
sccr_reg[464] = 8'h00;
sccr_reg[465] = 8'h00;
sccr_reg[466] = 8'h00;
sccr_reg[467] = 8'h00;
sccr_reg[468] = 8'h00;
sccr_reg[469] = 8'h00;
sccr_reg[470] = 8'h00;
sccr_reg[471] = 8'h00;
sccr_reg[472] = 8'h00;
sccr_reg[473] = 8'h00;
sccr_reg[474] = 8'h00;
sccr_reg[475] = 8'h00;
sccr_reg[476] = 8'h00;
sccr_reg[477] = 8'h00;
sccr_reg[478] = 8'h00;
sccr_reg[479] = 8'h00;
sccr_reg[480] = 8'h00;
sccr_reg[481] = 8'h00;
sccr_reg[482] = 8'h00;
sccr_reg[483] = 8'h00;
sccr_reg[484] = 8'h00;
sccr_reg[485] = 8'h00;
sccr_reg[486] = 8'h00;
sccr_reg[487] = 8'h00;
sccr_reg[488] = 8'h00;
sccr_reg[489] = 8'h00;
sccr_reg[490] = 8'h00;
sccr_reg[491] = 8'h00;
sccr_reg[492] = 8'h00;
sccr_reg[493] = 8'h00;
sccr_reg[494] = 8'h00;
sccr_reg[495] = 8'h00;
sccr_reg[496] = 8'h00;
sccr_reg[497] = 8'h00;
sccr_reg[498] = 8'h00;
sccr_reg[499] = 8'h00;
sccr_reg[500] = 8'h00;
sccr_reg[501] = 8'h00;
sccr_reg[502] = 8'h00;
sccr_reg[503] = 8'h00;
sccr_reg[504] = 8'h00;
sccr_reg[505] = 8'h00;
sccr_reg[506] = 8'h00;
sccr_reg[507] = 8'h00;
sccr_reg[508] = 8'h00;
sccr_reg[509] = 8'h00;
sccr_reg[510] = 8'h00;
sccr_reg[511] = 8'h00;
end